// q_sys_mSGDMA_0.v

// Generated using ACDS version 12.1sp1 243 at 2013.02.13.11:10:30

`timescale 1 ps / 1 ps
module q_sys_mSGDMA_0 (
		input  wire        reset_0_reset_n,                 //                  reset_0.reset_n
		output wire        dispatcher_write_csr_irq_irq,    // dispatcher_write_csr_irq.irq
		output wire [31:0] dma_read_master_address,         //          dma_read_master.address
		output wire        dma_read_master_read,            //                         .read
		output wire [7:0]  dma_read_master_byteenable,      //                         .byteenable
		input  wire [63:0] dma_read_master_readdata,        //                         .readdata
		input  wire        dma_read_master_waitrequest,     //                         .waitrequest
		input  wire        dma_read_master_readdatavalid,   //                         .readdatavalid
		output wire [5:0]  dma_read_master_burstcount,      //                         .burstcount
		output wire [31:0] dma_write_master_address,        //         dma_write_master.address
		output wire        dma_write_master_write,          //                         .write
		output wire [7:0]  dma_write_master_byteenable,     //                         .byteenable
		output wire [63:0] dma_write_master_writedata,      //                         .writedata
		input  wire        dma_write_master_waitrequest,    //                         .waitrequest
		output wire [5:0]  dma_write_master_burstcount,     //                         .burstcount
		output wire        mm_bridge_slv_waitrequest,       //            mm_bridge_slv.waitrequest
		output wire [31:0] mm_bridge_slv_readdata,          //                         .readdata
		output wire        mm_bridge_slv_readdatavalid,     //                         .readdatavalid
		input  wire [0:0]  mm_bridge_slv_burstcount,        //                         .burstcount
		input  wire [31:0] mm_bridge_slv_writedata,         //                         .writedata
		input  wire [19:0] mm_bridge_slv_address,           //                         .address
		input  wire        mm_bridge_slv_write,             //                         .write
		input  wire        mm_bridge_slv_read,              //                         .read
		input  wire [3:0]  mm_bridge_slv_byteenable,        //                         .byteenable
		input  wire        mm_bridge_slv_debugaccess,       //                         .debugaccess
		input  wire        reset_reset_n,                   //                    reset.reset_n
		output wire        reset_source_reset_n,            //             reset_source.reset_n
		input  wire        clk_clk,                         //                      clk.clk
		output wire        dispatcher_read_csr_irq_irq,     //  dispatcher_read_csr_irq.irq
		output wire        status_mon_out_cal_fail_mon,     //           status_mon_out.cal_fail_mon
		output wire        status_mon_out_cal_success_mon,  //                         .cal_success_mon
		output wire        status_mon_out_init_done_mon,    //                         .init_done_mon
		input  wire        clk_0_clk,                       //                    clk_0.clk
		input  wire        status_mon_in_local_init_done,   //            status_mon_in.local_init_done
		input  wire        status_mon_in_local_cal_success, //                         .local_cal_success
		input  wire        status_mon_in_local_cal_fail     //                         .local_cal_fail
	);

	wire          prbs_pattern_generator_st_pattern_output_valid;                                                         // prbs_pattern_generator:src_valid -> timing_adapter:in_valid
	wire   [63:0] prbs_pattern_generator_st_pattern_output_data;                                                          // prbs_pattern_generator:src_data -> timing_adapter:in_data
	wire          prbs_pattern_generator_st_pattern_output_ready;                                                         // timing_adapter:in_ready -> prbs_pattern_generator:src_ready
	wire          timing_adapter_out_valid;                                                                               // timing_adapter:out_valid -> dma_write_master:snk_valid
	wire   [63:0] timing_adapter_out_data;                                                                                // timing_adapter:out_data -> dma_write_master:snk_data
	wire          timing_adapter_out_ready;                                                                               // dma_write_master:snk_ready -> timing_adapter:out_ready
	wire          dispatcher_write_write_command_source_valid;                                                            // dispatcher_write:src_write_master_valid -> dma_write_master:snk_command_valid
	wire  [255:0] dispatcher_write_write_command_source_data;                                                             // dispatcher_write:src_write_master_data -> dma_write_master:snk_command_data
	wire          dispatcher_write_write_command_source_ready;                                                            // dma_write_master:snk_command_ready -> dispatcher_write:src_write_master_ready
	wire          dma_write_master_response_source_valid;                                                                 // dma_write_master:src_response_valid -> dispatcher_write:snk_write_master_valid
	wire  [255:0] dma_write_master_response_source_data;                                                                  // dma_write_master:src_response_data -> dispatcher_write:snk_write_master_data
	wire          dma_write_master_response_source_ready;                                                                 // dispatcher_write:snk_write_master_ready -> dma_write_master:src_response_ready
	wire          dma_read_master_data_source_valid;                                                                      // dma_read_master:src_valid -> prbs_pattern_checker:snk_valid
	wire   [63:0] dma_read_master_data_source_data;                                                                       // dma_read_master:src_data -> prbs_pattern_checker:snk_data
	wire          dma_read_master_data_source_ready;                                                                      // prbs_pattern_checker:snk_ready -> dma_read_master:src_ready
	wire          dispatcher_read_read_command_source_valid;                                                              // dispatcher_read:src_read_master_valid -> dma_read_master:snk_command_valid
	wire  [255:0] dispatcher_read_read_command_source_data;                                                               // dispatcher_read:src_read_master_data -> dma_read_master:snk_command_data
	wire          dispatcher_read_read_command_source_ready;                                                              // dma_read_master:snk_command_ready -> dispatcher_read:src_read_master_ready
	wire          dma_read_master_response_source_valid;                                                                  // dma_read_master:src_response_valid -> dispatcher_read:snk_read_master_valid
	wire  [255:0] dma_read_master_response_source_data;                                                                   // dma_read_master:src_response_data -> dispatcher_read:snk_read_master_data
	wire          dma_read_master_response_source_ready;                                                                  // dispatcher_read:snk_read_master_ready -> dma_read_master:src_response_ready
	wire    [0:0] mm_bridge_slv_m0_burstcount;                                                                            // mm_bridge_slv:m0_burstcount -> mm_bridge_slv_m0_translator:av_burstcount
	wire          mm_bridge_slv_m0_waitrequest;                                                                           // mm_bridge_slv_m0_translator:av_waitrequest -> mm_bridge_slv:m0_waitrequest
	wire   [19:0] mm_bridge_slv_m0_address;                                                                               // mm_bridge_slv:m0_address -> mm_bridge_slv_m0_translator:av_address
	wire   [31:0] mm_bridge_slv_m0_writedata;                                                                             // mm_bridge_slv:m0_writedata -> mm_bridge_slv_m0_translator:av_writedata
	wire          mm_bridge_slv_m0_write;                                                                                 // mm_bridge_slv:m0_write -> mm_bridge_slv_m0_translator:av_write
	wire          mm_bridge_slv_m0_read;                                                                                  // mm_bridge_slv:m0_read -> mm_bridge_slv_m0_translator:av_read
	wire   [31:0] mm_bridge_slv_m0_readdata;                                                                              // mm_bridge_slv_m0_translator:av_readdata -> mm_bridge_slv:m0_readdata
	wire          mm_bridge_slv_m0_debugaccess;                                                                           // mm_bridge_slv:m0_debugaccess -> mm_bridge_slv_m0_translator:av_debugaccess
	wire    [3:0] mm_bridge_slv_m0_byteenable;                                                                            // mm_bridge_slv:m0_byteenable -> mm_bridge_slv_m0_translator:av_byteenable
	wire          mm_bridge_slv_m0_readdatavalid;                                                                         // mm_bridge_slv_m0_translator:av_readdatavalid -> mm_bridge_slv:m0_readdatavalid
	wire   [31:0] prbs_pattern_generator_csr_translator_avalon_anti_slave_0_writedata;                                    // prbs_pattern_generator_csr_translator:av_writedata -> prbs_pattern_generator:csr_writedata
	wire    [2:0] prbs_pattern_generator_csr_translator_avalon_anti_slave_0_address;                                      // prbs_pattern_generator_csr_translator:av_address -> prbs_pattern_generator:csr_address
	wire          prbs_pattern_generator_csr_translator_avalon_anti_slave_0_write;                                        // prbs_pattern_generator_csr_translator:av_write -> prbs_pattern_generator:csr_write
	wire          prbs_pattern_generator_csr_translator_avalon_anti_slave_0_read;                                         // prbs_pattern_generator_csr_translator:av_read -> prbs_pattern_generator:csr_read
	wire   [31:0] prbs_pattern_generator_csr_translator_avalon_anti_slave_0_readdata;                                     // prbs_pattern_generator:csr_readdata -> prbs_pattern_generator_csr_translator:av_readdata
	wire    [3:0] prbs_pattern_generator_csr_translator_avalon_anti_slave_0_byteenable;                                   // prbs_pattern_generator_csr_translator:av_byteenable -> prbs_pattern_generator:csr_byteenable
	wire   [31:0] dispatcher_write_csr_translator_avalon_anti_slave_0_writedata;                                          // dispatcher_write_CSR_translator:av_writedata -> dispatcher_write:csr_writedata
	wire    [2:0] dispatcher_write_csr_translator_avalon_anti_slave_0_address;                                            // dispatcher_write_CSR_translator:av_address -> dispatcher_write:csr_address
	wire          dispatcher_write_csr_translator_avalon_anti_slave_0_write;                                              // dispatcher_write_CSR_translator:av_write -> dispatcher_write:csr_write
	wire          dispatcher_write_csr_translator_avalon_anti_slave_0_read;                                               // dispatcher_write_CSR_translator:av_read -> dispatcher_write:csr_read
	wire   [31:0] dispatcher_write_csr_translator_avalon_anti_slave_0_readdata;                                           // dispatcher_write:csr_readdata -> dispatcher_write_CSR_translator:av_readdata
	wire    [3:0] dispatcher_write_csr_translator_avalon_anti_slave_0_byteenable;                                         // dispatcher_write_CSR_translator:av_byteenable -> dispatcher_write:csr_byteenable
	wire          dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_waitrequest;                           // dispatcher_write:descriptor_waitrequest -> dispatcher_write_Descriptor_Slave_translator:av_waitrequest
	wire  [127:0] dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_writedata;                             // dispatcher_write_Descriptor_Slave_translator:av_writedata -> dispatcher_write:descriptor_writedata
	wire          dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_write;                                 // dispatcher_write_Descriptor_Slave_translator:av_write -> dispatcher_write:descriptor_write
	wire   [15:0] dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_byteenable;                            // dispatcher_write_Descriptor_Slave_translator:av_byteenable -> dispatcher_write:descriptor_byteenable
	wire   [31:0] prbs_pattern_checker_csr_translator_avalon_anti_slave_0_writedata;                                      // prbs_pattern_checker_csr_translator:av_writedata -> prbs_pattern_checker:csr_writedata
	wire    [3:0] prbs_pattern_checker_csr_translator_avalon_anti_slave_0_address;                                        // prbs_pattern_checker_csr_translator:av_address -> prbs_pattern_checker:csr_address
	wire          prbs_pattern_checker_csr_translator_avalon_anti_slave_0_write;                                          // prbs_pattern_checker_csr_translator:av_write -> prbs_pattern_checker:csr_write
	wire          prbs_pattern_checker_csr_translator_avalon_anti_slave_0_read;                                           // prbs_pattern_checker_csr_translator:av_read -> prbs_pattern_checker:csr_read
	wire   [31:0] prbs_pattern_checker_csr_translator_avalon_anti_slave_0_readdata;                                       // prbs_pattern_checker:csr_readdata -> prbs_pattern_checker_csr_translator:av_readdata
	wire    [3:0] prbs_pattern_checker_csr_translator_avalon_anti_slave_0_byteenable;                                     // prbs_pattern_checker_csr_translator:av_byteenable -> prbs_pattern_checker:csr_byteenable
	wire   [31:0] dispatcher_read_csr_translator_avalon_anti_slave_0_writedata;                                           // dispatcher_read_CSR_translator:av_writedata -> dispatcher_read:csr_writedata
	wire    [2:0] dispatcher_read_csr_translator_avalon_anti_slave_0_address;                                             // dispatcher_read_CSR_translator:av_address -> dispatcher_read:csr_address
	wire          dispatcher_read_csr_translator_avalon_anti_slave_0_write;                                               // dispatcher_read_CSR_translator:av_write -> dispatcher_read:csr_write
	wire          dispatcher_read_csr_translator_avalon_anti_slave_0_read;                                                // dispatcher_read_CSR_translator:av_read -> dispatcher_read:csr_read
	wire   [31:0] dispatcher_read_csr_translator_avalon_anti_slave_0_readdata;                                            // dispatcher_read:csr_readdata -> dispatcher_read_CSR_translator:av_readdata
	wire    [3:0] dispatcher_read_csr_translator_avalon_anti_slave_0_byteenable;                                          // dispatcher_read_CSR_translator:av_byteenable -> dispatcher_read:csr_byteenable
	wire          dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_waitrequest;                            // dispatcher_read:descriptor_waitrequest -> dispatcher_read_Descriptor_Slave_translator:av_waitrequest
	wire  [127:0] dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_writedata;                              // dispatcher_read_Descriptor_Slave_translator:av_writedata -> dispatcher_read:descriptor_writedata
	wire          dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_write;                                  // dispatcher_read_Descriptor_Slave_translator:av_write -> dispatcher_read:descriptor_write
	wire   [15:0] dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_byteenable;                             // dispatcher_read_Descriptor_Slave_translator:av_byteenable -> dispatcher_read:descriptor_byteenable
	wire   [31:0] status_mon_0_slv_translator_avalon_anti_slave_0_writedata;                                              // status_mon_0_slv_translator:av_writedata -> status_mon_0:slv_data_write
	wire    [1:0] status_mon_0_slv_translator_avalon_anti_slave_0_address;                                                // status_mon_0_slv_translator:av_address -> status_mon_0:slv_address
	wire          status_mon_0_slv_translator_avalon_anti_slave_0_chipselect;                                             // status_mon_0_slv_translator:av_chipselect -> status_mon_0:slv_cs_n
	wire          status_mon_0_slv_translator_avalon_anti_slave_0_write;                                                  // status_mon_0_slv_translator:av_write -> status_mon_0:slv_write_n
	wire          status_mon_0_slv_translator_avalon_anti_slave_0_read;                                                   // status_mon_0_slv_translator:av_read -> status_mon_0:slv_read_n
	wire   [31:0] status_mon_0_slv_translator_avalon_anti_slave_0_readdata;                                               // status_mon_0:slv_data_read -> status_mon_0_slv_translator:av_readdata
	wire          frequency_counter_0_csr_translator_avalon_anti_slave_0_waitrequest;                                     // frequency_counter_0:csr_waitrequest -> frequency_counter_0_csr_translator:av_waitrequest
	wire    [3:0] frequency_counter_0_csr_translator_avalon_anti_slave_0_address;                                         // frequency_counter_0_csr_translator:av_address -> frequency_counter_0:csr_address
	wire          frequency_counter_0_csr_translator_avalon_anti_slave_0_read;                                            // frequency_counter_0_csr_translator:av_read -> frequency_counter_0:csr_read
	wire   [31:0] frequency_counter_0_csr_translator_avalon_anti_slave_0_readdata;                                        // frequency_counter_0:csr_readdata -> frequency_counter_0_csr_translator:av_readdata
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire    [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_0_s1_translator:av_address -> timer_0:address
	wire          timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire          timer_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_0_s1_translator:av_write -> timer_0:write_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_waitrequest;                                      // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_bridge_slv_m0_translator:uav_waitrequest
	wire    [2:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_burstcount;                                       // mm_bridge_slv_m0_translator:uav_burstcount -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_writedata;                                        // mm_bridge_slv_m0_translator:uav_writedata -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [19:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_address;                                          // mm_bridge_slv_m0_translator:uav_address -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_address
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_lock;                                             // mm_bridge_slv_m0_translator:uav_lock -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_write;                                            // mm_bridge_slv_m0_translator:uav_write -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_write
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_read;                                             // mm_bridge_slv_m0_translator:uav_read -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_readdata;                                         // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_bridge_slv_m0_translator:uav_readdata
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_debugaccess;                                      // mm_bridge_slv_m0_translator:uav_debugaccess -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_byteenable;                                       // mm_bridge_slv_m0_translator:uav_byteenable -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_readdatavalid;                                    // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_bridge_slv_m0_translator:uav_readdatavalid
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // prbs_pattern_generator_csr_translator:uav_waitrequest -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> prbs_pattern_generator_csr_translator:uav_burstcount
	wire   [31:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                      // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> prbs_pattern_generator_csr_translator:uav_writedata
	wire   [19:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_address;                        // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_address -> prbs_pattern_generator_csr_translator:uav_address
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_write;                          // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_write -> prbs_pattern_generator_csr_translator:uav_write
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_lock;                           // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_lock -> prbs_pattern_generator_csr_translator:uav_lock
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_read;                           // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_read -> prbs_pattern_generator_csr_translator:uav_read
	wire   [31:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                       // prbs_pattern_generator_csr_translator:uav_readdata -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // prbs_pattern_generator_csr_translator:uav_readdatavalid -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prbs_pattern_generator_csr_translator:uav_debugaccess
	wire    [3:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> prbs_pattern_generator_csr_translator:uav_byteenable
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                    // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // dispatcher_write_CSR_translator:uav_waitrequest -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_burstcount -> dispatcher_write_CSR_translator:uav_burstcount
	wire   [31:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                            // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_writedata -> dispatcher_write_CSR_translator:uav_writedata
	wire   [19:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_address;                              // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_address -> dispatcher_write_CSR_translator:uav_address
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_write;                                // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_write -> dispatcher_write_CSR_translator:uav_write
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                 // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_lock -> dispatcher_write_CSR_translator:uav_lock
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_read;                                 // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_read -> dispatcher_write_CSR_translator:uav_read
	wire   [31:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                             // dispatcher_write_CSR_translator:uav_readdata -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // dispatcher_write_CSR_translator:uav_readdatavalid -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dispatcher_write_CSR_translator:uav_debugaccess
	wire    [3:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:m0_byteenable -> dispatcher_write_CSR_translator:uav_byteenable
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_source_valid -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                          // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_source_data -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // dispatcher_write_Descriptor_Slave_translator:uav_waitrequest -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [4:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dispatcher_write_Descriptor_Slave_translator:uav_burstcount
	wire  [127:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dispatcher_write_Descriptor_Slave_translator:uav_writedata
	wire   [19:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_address -> dispatcher_write_Descriptor_Slave_translator:uav_address
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_write -> dispatcher_write_Descriptor_Slave_translator:uav_write
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_lock -> dispatcher_write_Descriptor_Slave_translator:uav_lock
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_read -> dispatcher_write_Descriptor_Slave_translator:uav_read
	wire  [127:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // dispatcher_write_Descriptor_Slave_translator:uav_readdata -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // dispatcher_write_Descriptor_Slave_translator:uav_readdatavalid -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dispatcher_write_Descriptor_Slave_translator:uav_debugaccess
	wire   [15:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dispatcher_write_Descriptor_Slave_translator:uav_byteenable
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [207:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [207:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [127:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // prbs_pattern_checker_csr_translator:uav_waitrequest -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> prbs_pattern_checker_csr_translator:uav_burstcount
	wire   [31:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                        // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> prbs_pattern_checker_csr_translator:uav_writedata
	wire   [19:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_address;                          // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_address -> prbs_pattern_checker_csr_translator:uav_address
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_write;                            // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_write -> prbs_pattern_checker_csr_translator:uav_write
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_lock;                             // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_lock -> prbs_pattern_checker_csr_translator:uav_lock
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_read;                             // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_read -> prbs_pattern_checker_csr_translator:uav_read
	wire   [31:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                         // prbs_pattern_checker_csr_translator:uav_readdata -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // prbs_pattern_checker_csr_translator:uav_readdatavalid -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prbs_pattern_checker_csr_translator:uav_debugaccess
	wire    [3:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> prbs_pattern_checker_csr_translator:uav_byteenable
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                      // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // dispatcher_read_CSR_translator:uav_waitrequest -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_burstcount -> dispatcher_read_CSR_translator:uav_burstcount
	wire   [31:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                             // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_writedata -> dispatcher_read_CSR_translator:uav_writedata
	wire   [19:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_address;                               // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_address -> dispatcher_read_CSR_translator:uav_address
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_write;                                 // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_write -> dispatcher_read_CSR_translator:uav_write
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                  // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_lock -> dispatcher_read_CSR_translator:uav_lock
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_read;                                  // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_read -> dispatcher_read_CSR_translator:uav_read
	wire   [31:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                              // dispatcher_read_CSR_translator:uav_readdata -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // dispatcher_read_CSR_translator:uav_readdatavalid -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dispatcher_read_CSR_translator:uav_debugaccess
	wire    [3:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:m0_byteenable -> dispatcher_read_CSR_translator:uav_byteenable
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_source_valid -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                           // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_source_data -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // dispatcher_read_Descriptor_Slave_translator:uav_waitrequest -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [4:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dispatcher_read_Descriptor_Slave_translator:uav_burstcount
	wire  [127:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dispatcher_read_Descriptor_Slave_translator:uav_writedata
	wire   [19:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_address -> dispatcher_read_Descriptor_Slave_translator:uav_address
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_write -> dispatcher_read_Descriptor_Slave_translator:uav_write
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_lock -> dispatcher_read_Descriptor_Slave_translator:uav_lock
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_read -> dispatcher_read_Descriptor_Slave_translator:uav_read
	wire  [127:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // dispatcher_read_Descriptor_Slave_translator:uav_readdata -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // dispatcher_read_Descriptor_Slave_translator:uav_readdatavalid -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dispatcher_read_Descriptor_Slave_translator:uav_debugaccess
	wire   [15:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dispatcher_read_Descriptor_Slave_translator:uav_byteenable
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [207:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [207:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [127:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // status_mon_0_slv_translator:uav_waitrequest -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_burstcount -> status_mon_0_slv_translator:uav_burstcount
	wire   [31:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_writedata;                                // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_writedata -> status_mon_0_slv_translator:uav_writedata
	wire   [19:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_address;                                  // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_address -> status_mon_0_slv_translator:uav_address
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_write;                                    // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_write -> status_mon_0_slv_translator:uav_write
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_lock;                                     // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_lock -> status_mon_0_slv_translator:uav_lock
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_read;                                     // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_read -> status_mon_0_slv_translator:uav_read
	wire   [31:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // status_mon_0_slv_translator:uav_readdata -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // status_mon_0_slv_translator:uav_readdatavalid -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_debugaccess -> status_mon_0_slv_translator:uav_debugaccess
	wire    [3:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // status_mon_0_slv_translator_avalon_universal_slave_0_agent:m0_byteenable -> status_mon_0_slv_translator:uav_byteenable
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_source_valid -> status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_data;                              // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_source_data -> status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rf_sink_ready -> status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // frequency_counter_0_csr_translator:uav_waitrequest -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> frequency_counter_0_csr_translator:uav_burstcount
	wire   [31:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                         // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> frequency_counter_0_csr_translator:uav_writedata
	wire   [19:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_address;                           // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_address -> frequency_counter_0_csr_translator:uav_address
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_write;                             // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_write -> frequency_counter_0_csr_translator:uav_write
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_lock;                              // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_lock -> frequency_counter_0_csr_translator:uav_lock
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_read;                              // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_read -> frequency_counter_0_csr_translator:uav_read
	wire   [31:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                          // frequency_counter_0_csr_translator:uav_readdata -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // frequency_counter_0_csr_translator:uav_readdatavalid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> frequency_counter_0_csr_translator:uav_debugaccess
	wire    [3:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> frequency_counter_0_csr_translator:uav_byteenable
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                       // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire   [19:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire    [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_valid;                                   // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [98:0] mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_data;                                    // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router:sink_ready -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [98:0] addr_router_src_data;                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire    [8:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [98:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [8:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                  // mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> [addr_router:reset, agent_pipeline:reset, agent_pipeline_001:reset, agent_pipeline_002:reset, agent_pipeline_003:reset, agent_pipeline_004:reset, agent_pipeline_005:reset, agent_pipeline_006:reset, agent_pipeline_007:reset, agent_pipeline_008:reset, agent_pipeline_009:reset, agent_pipeline_010:reset, agent_pipeline_011:reset, agent_pipeline_012:reset, agent_pipeline_013:reset, cmd_xbar_demux:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, dispatcher_read:reset, dispatcher_read_CSR_translator:reset, dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:reset, dispatcher_read_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dispatcher_read_Descriptor_Slave_translator:reset, dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:reset, dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dispatcher_write:reset, dispatcher_write_CSR_translator:reset, dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:reset, dispatcher_write_CSR_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dispatcher_write_Descriptor_Slave_translator:reset, dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:reset, dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_read_master:reset, dma_write_master:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, limiter:reset, limiter_pipeline:reset, limiter_pipeline_001:reset, mm_bridge_slv:reset, mm_bridge_slv_m0_translator:reset, mm_bridge_slv_m0_translator_avalon_universal_master_0_agent:reset, mux_pipeline:reset, mux_pipeline_001:reset, mux_pipeline_002:reset, mux_pipeline_003:reset, mux_pipeline_004:reset, mux_pipeline_005:reset, mux_pipeline_006:reset, mux_pipeline_009:reset, mux_pipeline_010:reset, mux_pipeline_011:reset, mux_pipeline_012:reset, mux_pipeline_013:reset, mux_pipeline_014:reset, mux_pipeline_015:reset, mux_pipeline_016:reset, mux_pipeline_017:reset, prbs_pattern_checker:reset, prbs_pattern_checker_csr_translator:reset, prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:reset, prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prbs_pattern_generator:reset, prbs_pattern_generator_csr_translator:reset, prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:reset, prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset, status_mon_0:slv_reset_n, status_mon_0_slv_translator:reset, status_mon_0_slv_translator_avalon_universal_slave_0_agent:reset, status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timing_adapter:reset_n, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_001_reset_out_reset;                                                                     // rst_controller_001:reset_out -> [agent_pipeline_014:reset, agent_pipeline_015:reset, crosser:out_reset, crosser_002:in_reset, frequency_counter_0:reset_n, frequency_counter_0_csr_translator:reset, frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:reset, frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, mux_pipeline_007:reset, rsp_xbar_demux_007:reset]
	wire          rst_controller_002_reset_out_reset;                                                                     // rst_controller_002:reset_out -> frequency_counter_0:sample_reset_n
	wire          rst_controller_003_reset_out_reset;                                                                     // rst_controller_003:reset_out -> [agent_pipeline_016:reset, agent_pipeline_017:reset, crosser_001:out_reset, crosser_003:in_reset, id_router_008:reset, mux_pipeline_008:reset, rsp_xbar_demux_008:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [98:0] id_router_src_data;                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [8:0] id_router_src_channel;                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [98:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [8:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [98:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [8:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [98:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [8:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          id_router_006_src_endofpacket;                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [98:0] id_router_006_src_data;                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [8:0] id_router_006_src_channel;                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          id_router_007_src_endofpacket;                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [98:0] id_router_007_src_data;                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [8:0] id_router_007_src_channel;                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          id_router_008_src_endofpacket;                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [98:0] id_router_008_src_data;                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [8:0] id_router_008_src_channel;                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          mux_pipeline_002_source0_ready;                                                                         // width_adapter:in_ready -> mux_pipeline_002:out_ready
	wire          id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_002_src_valid;                                                                                // id_router_002:src_valid -> width_adapter_001:in_valid
	wire          id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [206:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> width_adapter_001:in_data
	wire    [8:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> width_adapter_001:in_channel
	wire          id_router_002_src_ready;                                                                                // width_adapter_001:in_ready -> id_router_002:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [98:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_001_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire    [8:0] width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          mux_pipeline_005_source0_ready;                                                                         // width_adapter_002:in_ready -> mux_pipeline_005:out_ready
	wire          id_router_005_src_endofpacket;                                                                          // id_router_005:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_005_src_valid;                                                                                // id_router_005:src_valid -> width_adapter_003:in_valid
	wire          id_router_005_src_startofpacket;                                                                        // id_router_005:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [206:0] id_router_005_src_data;                                                                                 // id_router_005:src_data -> width_adapter_003:in_data
	wire    [8:0] id_router_005_src_channel;                                                                              // id_router_005:src_channel -> width_adapter_003:in_channel
	wire          id_router_005_src_ready;                                                                                // width_adapter_003:in_ready -> id_router_005:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> rsp_xbar_demux_005:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [98:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> rsp_xbar_demux_005:sink_data
	wire          width_adapter_003_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> width_adapter_003:out_ready
	wire    [8:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> rsp_xbar_demux_005:sink_channel
	wire          cmd_xbar_demux_src7_endofpacket;                                                                        // cmd_xbar_demux:src7_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                              // cmd_xbar_demux:src7_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                      // cmd_xbar_demux:src7_startofpacket -> crosser:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src7_data;                                                                               // cmd_xbar_demux:src7_data -> crosser:in_data
	wire    [8:0] cmd_xbar_demux_src7_channel;                                                                            // cmd_xbar_demux:src7_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src7_ready;                                                                              // crosser:in_ready -> cmd_xbar_demux:src7_ready
	wire          cmd_xbar_demux_src8_endofpacket;                                                                        // cmd_xbar_demux:src8_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                              // cmd_xbar_demux:src8_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                      // cmd_xbar_demux:src8_startofpacket -> crosser_001:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src8_data;                                                                               // cmd_xbar_demux:src8_data -> crosser_001:in_data
	wire    [8:0] cmd_xbar_demux_src8_channel;                                                                            // cmd_xbar_demux:src8_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_src8_ready;                                                                              // crosser_001:in_ready -> cmd_xbar_demux:src8_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                    // rsp_xbar_demux_007:src0_endofpacket -> crosser_002:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                          // rsp_xbar_demux_007:src0_valid -> crosser_002:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                  // rsp_xbar_demux_007:src0_startofpacket -> crosser_002:in_startofpacket
	wire   [98:0] rsp_xbar_demux_007_src0_data;                                                                           // rsp_xbar_demux_007:src0_data -> crosser_002:in_data
	wire    [8:0] rsp_xbar_demux_007_src0_channel;                                                                        // rsp_xbar_demux_007:src0_channel -> crosser_002:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                          // crosser_002:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                    // rsp_xbar_demux_008:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                          // rsp_xbar_demux_008:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                  // rsp_xbar_demux_008:src0_startofpacket -> crosser_003:in_startofpacket
	wire   [98:0] rsp_xbar_demux_008_src0_data;                                                                           // rsp_xbar_demux_008:src0_data -> crosser_003:in_data
	wire    [8:0] rsp_xbar_demux_008_src0_channel;                                                                        // rsp_xbar_demux_008:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                          // crosser_003:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          limiter_pipeline_source0_endofpacket;                                                                   // limiter_pipeline:out_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_pipeline_source0_valid;                                                                         // limiter_pipeline:out_valid -> cmd_xbar_demux:sink_valid
	wire          limiter_pipeline_source0_startofpacket;                                                                 // limiter_pipeline:out_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [98:0] limiter_pipeline_source0_data;                                                                          // limiter_pipeline:out_data -> cmd_xbar_demux:sink_data
	wire    [8:0] limiter_pipeline_source0_channel;                                                                       // limiter_pipeline:out_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_pipeline_source0_ready;                                                                         // cmd_xbar_demux:sink_ready -> limiter_pipeline:out_ready
	wire          limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> limiter_pipeline:in_endofpacket
	wire    [0:0] limiter_cmd_src_valid;                                                                                  // limiter:cmd_src_valid -> limiter_pipeline:in_valid
	wire          limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> limiter_pipeline:in_startofpacket
	wire   [98:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> limiter_pipeline:in_data
	wire    [8:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> limiter_pipeline:in_channel
	wire          limiter_cmd_src_ready;                                                                                  // limiter_pipeline:in_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                           // rsp_xbar_mux:src_endofpacket -> limiter_pipeline_001:in_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                 // rsp_xbar_mux:src_valid -> limiter_pipeline_001:in_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                         // rsp_xbar_mux:src_startofpacket -> limiter_pipeline_001:in_startofpacket
	wire   [98:0] rsp_xbar_mux_src_data;                                                                                  // rsp_xbar_mux:src_data -> limiter_pipeline_001:in_data
	wire    [8:0] rsp_xbar_mux_src_channel;                                                                               // rsp_xbar_mux:src_channel -> limiter_pipeline_001:in_channel
	wire          rsp_xbar_mux_src_ready;                                                                                 // limiter_pipeline_001:in_ready -> rsp_xbar_mux:src_ready
	wire          limiter_pipeline_001_source0_endofpacket;                                                               // limiter_pipeline_001:out_endofpacket -> limiter:rsp_sink_endofpacket
	wire          limiter_pipeline_001_source0_valid;                                                                     // limiter_pipeline_001:out_valid -> limiter:rsp_sink_valid
	wire          limiter_pipeline_001_source0_startofpacket;                                                             // limiter_pipeline_001:out_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [98:0] limiter_pipeline_001_source0_data;                                                                      // limiter_pipeline_001:out_data -> limiter:rsp_sink_data
	wire    [8:0] limiter_pipeline_001_source0_channel;                                                                   // limiter_pipeline_001:out_channel -> limiter:rsp_sink_channel
	wire          limiter_pipeline_001_source0_ready;                                                                     // limiter:rsp_sink_ready -> limiter_pipeline_001:out_ready
	wire          mux_pipeline_source0_ready;                                                                             // agent_pipeline:in_ready -> mux_pipeline:out_ready
	wire          agent_pipeline_source0_endofpacket;                                                                     // agent_pipeline:out_endofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_source0_valid;                                                                           // agent_pipeline:out_valid -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_source0_startofpacket;                                                                   // agent_pipeline:out_startofpacket -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_source0_data;                                                                            // agent_pipeline:out_data -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_source0_channel;                                                                         // agent_pipeline:out_channel -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_source0_ready;                                                                           // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline:out_ready
	wire          agent_pipeline_001_source0_endofpacket;                                                                 // agent_pipeline_001:out_endofpacket -> id_router:sink_endofpacket
	wire          agent_pipeline_001_source0_valid;                                                                       // agent_pipeline_001:out_valid -> id_router:sink_valid
	wire          agent_pipeline_001_source0_startofpacket;                                                               // agent_pipeline_001:out_startofpacket -> id_router:sink_startofpacket
	wire   [98:0] agent_pipeline_001_source0_data;                                                                        // agent_pipeline_001:out_data -> id_router:sink_data
	wire          agent_pipeline_001_source0_ready;                                                                       // id_router:sink_ready -> agent_pipeline_001:out_ready
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_001:in_endofpacket
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_valid;                          // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_001:in_valid
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_001:in_startofpacket
	wire   [98:0] prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_data;                           // prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_001:in_data
	wire          prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_ready;                          // agent_pipeline_001:in_ready -> prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_001_source0_ready;                                                                         // agent_pipeline_002:in_ready -> mux_pipeline_001:out_ready
	wire          agent_pipeline_002_source0_endofpacket;                                                                 // agent_pipeline_002:out_endofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_002_source0_valid;                                                                       // agent_pipeline_002:out_valid -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_002_source0_startofpacket;                                                               // agent_pipeline_002:out_startofpacket -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_002_source0_data;                                                                        // agent_pipeline_002:out_data -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_002_source0_channel;                                                                     // agent_pipeline_002:out_channel -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_002_source0_ready;                                                                       // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_002:out_ready
	wire          agent_pipeline_003_source0_endofpacket;                                                                 // agent_pipeline_003:out_endofpacket -> id_router_001:sink_endofpacket
	wire          agent_pipeline_003_source0_valid;                                                                       // agent_pipeline_003:out_valid -> id_router_001:sink_valid
	wire          agent_pipeline_003_source0_startofpacket;                                                               // agent_pipeline_003:out_startofpacket -> id_router_001:sink_startofpacket
	wire   [98:0] agent_pipeline_003_source0_data;                                                                        // agent_pipeline_003:out_data -> id_router_001:sink_data
	wire          agent_pipeline_003_source0_ready;                                                                       // id_router_001:sink_ready -> agent_pipeline_003:out_ready
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_003:in_endofpacket
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_003:in_valid
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_003:in_startofpacket
	wire   [98:0] dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_data;                                 // dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_003:in_data
	wire          dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                // agent_pipeline_003:in_ready -> dispatcher_write_CSR_translator_avalon_universal_slave_0_agent:rp_ready
	wire          width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> agent_pipeline_004:in_endofpacket
	wire          width_adapter_src_valid;                                                                                // width_adapter:out_valid -> agent_pipeline_004:in_valid
	wire          width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> agent_pipeline_004:in_startofpacket
	wire  [206:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> agent_pipeline_004:in_data
	wire          width_adapter_src_ready;                                                                                // agent_pipeline_004:in_ready -> width_adapter:out_ready
	wire    [8:0] width_adapter_src_channel;                                                                              // width_adapter:out_channel -> agent_pipeline_004:in_channel
	wire          agent_pipeline_004_source0_endofpacket;                                                                 // agent_pipeline_004:out_endofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_004_source0_valid;                                                                       // agent_pipeline_004:out_valid -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_004_source0_startofpacket;                                                               // agent_pipeline_004:out_startofpacket -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [206:0] agent_pipeline_004_source0_data;                                                                        // agent_pipeline_004:out_data -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_004_source0_channel;                                                                     // agent_pipeline_004:out_channel -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_004_source0_ready;                                                                       // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_004:out_ready
	wire          agent_pipeline_005_source0_endofpacket;                                                                 // agent_pipeline_005:out_endofpacket -> id_router_002:sink_endofpacket
	wire          agent_pipeline_005_source0_valid;                                                                       // agent_pipeline_005:out_valid -> id_router_002:sink_valid
	wire          agent_pipeline_005_source0_startofpacket;                                                               // agent_pipeline_005:out_startofpacket -> id_router_002:sink_startofpacket
	wire  [206:0] agent_pipeline_005_source0_data;                                                                        // agent_pipeline_005:out_data -> id_router_002:sink_data
	wire          agent_pipeline_005_source0_ready;                                                                       // id_router_002:sink_ready -> agent_pipeline_005:out_ready
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_005:in_endofpacket
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_005:in_valid
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_005:in_startofpacket
	wire  [206:0] dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_005:in_data
	wire          dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // agent_pipeline_005:in_ready -> dispatcher_write_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_003_source0_ready;                                                                         // agent_pipeline_006:in_ready -> mux_pipeline_003:out_ready
	wire          agent_pipeline_006_source0_endofpacket;                                                                 // agent_pipeline_006:out_endofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_006_source0_valid;                                                                       // agent_pipeline_006:out_valid -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_006_source0_startofpacket;                                                               // agent_pipeline_006:out_startofpacket -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_006_source0_data;                                                                        // agent_pipeline_006:out_data -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_006_source0_channel;                                                                     // agent_pipeline_006:out_channel -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_006_source0_ready;                                                                       // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_006:out_ready
	wire          agent_pipeline_007_source0_endofpacket;                                                                 // agent_pipeline_007:out_endofpacket -> id_router_003:sink_endofpacket
	wire          agent_pipeline_007_source0_valid;                                                                       // agent_pipeline_007:out_valid -> id_router_003:sink_valid
	wire          agent_pipeline_007_source0_startofpacket;                                                               // agent_pipeline_007:out_startofpacket -> id_router_003:sink_startofpacket
	wire   [98:0] agent_pipeline_007_source0_data;                                                                        // agent_pipeline_007:out_data -> id_router_003:sink_data
	wire          agent_pipeline_007_source0_ready;                                                                       // id_router_003:sink_ready -> agent_pipeline_007:out_ready
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_007:in_endofpacket
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_valid;                            // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_007:in_valid
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_007:in_startofpacket
	wire   [98:0] prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_data;                             // prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_007:in_data
	wire          prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_ready;                            // agent_pipeline_007:in_ready -> prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_004_source0_ready;                                                                         // agent_pipeline_008:in_ready -> mux_pipeline_004:out_ready
	wire          agent_pipeline_008_source0_endofpacket;                                                                 // agent_pipeline_008:out_endofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_008_source0_valid;                                                                       // agent_pipeline_008:out_valid -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_008_source0_startofpacket;                                                               // agent_pipeline_008:out_startofpacket -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_008_source0_data;                                                                        // agent_pipeline_008:out_data -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_008_source0_channel;                                                                     // agent_pipeline_008:out_channel -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_008_source0_ready;                                                                       // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_008:out_ready
	wire          agent_pipeline_009_source0_endofpacket;                                                                 // agent_pipeline_009:out_endofpacket -> id_router_004:sink_endofpacket
	wire          agent_pipeline_009_source0_valid;                                                                       // agent_pipeline_009:out_valid -> id_router_004:sink_valid
	wire          agent_pipeline_009_source0_startofpacket;                                                               // agent_pipeline_009:out_startofpacket -> id_router_004:sink_startofpacket
	wire   [98:0] agent_pipeline_009_source0_data;                                                                        // agent_pipeline_009:out_data -> id_router_004:sink_data
	wire          agent_pipeline_009_source0_ready;                                                                       // id_router_004:sink_ready -> agent_pipeline_009:out_ready
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_009:in_endofpacket
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                 // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_009:in_valid
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_009:in_startofpacket
	wire   [98:0] dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_data;                                  // dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_009:in_data
	wire          dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                 // agent_pipeline_009:in_ready -> dispatcher_read_CSR_translator_avalon_universal_slave_0_agent:rp_ready
	wire          width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> agent_pipeline_010:in_endofpacket
	wire          width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> agent_pipeline_010:in_valid
	wire          width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> agent_pipeline_010:in_startofpacket
	wire  [206:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> agent_pipeline_010:in_data
	wire          width_adapter_002_src_ready;                                                                            // agent_pipeline_010:in_ready -> width_adapter_002:out_ready
	wire    [8:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> agent_pipeline_010:in_channel
	wire          agent_pipeline_010_source0_endofpacket;                                                                 // agent_pipeline_010:out_endofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_010_source0_valid;                                                                       // agent_pipeline_010:out_valid -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_010_source0_startofpacket;                                                               // agent_pipeline_010:out_startofpacket -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [206:0] agent_pipeline_010_source0_data;                                                                        // agent_pipeline_010:out_data -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_010_source0_channel;                                                                     // agent_pipeline_010:out_channel -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_010_source0_ready;                                                                       // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_010:out_ready
	wire          agent_pipeline_011_source0_endofpacket;                                                                 // agent_pipeline_011:out_endofpacket -> id_router_005:sink_endofpacket
	wire          agent_pipeline_011_source0_valid;                                                                       // agent_pipeline_011:out_valid -> id_router_005:sink_valid
	wire          agent_pipeline_011_source0_startofpacket;                                                               // agent_pipeline_011:out_startofpacket -> id_router_005:sink_startofpacket
	wire  [206:0] agent_pipeline_011_source0_data;                                                                        // agent_pipeline_011:out_data -> id_router_005:sink_data
	wire          agent_pipeline_011_source0_ready;                                                                       // id_router_005:sink_ready -> agent_pipeline_011:out_ready
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_011:in_endofpacket
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_011:in_valid
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_011:in_startofpacket
	wire  [206:0] dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_011:in_data
	wire          dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // agent_pipeline_011:in_ready -> dispatcher_read_Descriptor_Slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_006_source0_ready;                                                                         // agent_pipeline_012:in_ready -> mux_pipeline_006:out_ready
	wire          agent_pipeline_012_source0_endofpacket;                                                                 // agent_pipeline_012:out_endofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_012_source0_valid;                                                                       // agent_pipeline_012:out_valid -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_012_source0_startofpacket;                                                               // agent_pipeline_012:out_startofpacket -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_012_source0_data;                                                                        // agent_pipeline_012:out_data -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_012_source0_channel;                                                                     // agent_pipeline_012:out_channel -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_012_source0_ready;                                                                       // status_mon_0_slv_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_012:out_ready
	wire          agent_pipeline_013_source0_endofpacket;                                                                 // agent_pipeline_013:out_endofpacket -> id_router_006:sink_endofpacket
	wire          agent_pipeline_013_source0_valid;                                                                       // agent_pipeline_013:out_valid -> id_router_006:sink_valid
	wire          agent_pipeline_013_source0_startofpacket;                                                               // agent_pipeline_013:out_startofpacket -> id_router_006:sink_startofpacket
	wire   [98:0] agent_pipeline_013_source0_data;                                                                        // agent_pipeline_013:out_data -> id_router_006:sink_data
	wire          agent_pipeline_013_source0_ready;                                                                       // id_router_006:sink_ready -> agent_pipeline_013:out_ready
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_013:in_endofpacket
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_valid;                                    // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_013:in_valid
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_013:in_startofpacket
	wire   [98:0] status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_data;                                     // status_mon_0_slv_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_013:in_data
	wire          status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_ready;                                    // agent_pipeline_013:in_ready -> status_mon_0_slv_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_007_source0_ready;                                                                         // agent_pipeline_014:in_ready -> mux_pipeline_007:out_ready
	wire          agent_pipeline_014_source0_endofpacket;                                                                 // agent_pipeline_014:out_endofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_014_source0_valid;                                                                       // agent_pipeline_014:out_valid -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_014_source0_startofpacket;                                                               // agent_pipeline_014:out_startofpacket -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_014_source0_data;                                                                        // agent_pipeline_014:out_data -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_014_source0_channel;                                                                     // agent_pipeline_014:out_channel -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_014_source0_ready;                                                                       // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_014:out_ready
	wire          agent_pipeline_015_source0_endofpacket;                                                                 // agent_pipeline_015:out_endofpacket -> id_router_007:sink_endofpacket
	wire          agent_pipeline_015_source0_valid;                                                                       // agent_pipeline_015:out_valid -> id_router_007:sink_valid
	wire          agent_pipeline_015_source0_startofpacket;                                                               // agent_pipeline_015:out_startofpacket -> id_router_007:sink_startofpacket
	wire   [98:0] agent_pipeline_015_source0_data;                                                                        // agent_pipeline_015:out_data -> id_router_007:sink_data
	wire          agent_pipeline_015_source0_ready;                                                                       // id_router_007:sink_ready -> agent_pipeline_015:out_ready
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_015:in_endofpacket
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_valid;                             // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_015:in_valid
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_015:in_startofpacket
	wire   [98:0] frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_data;                              // frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_015:in_data
	wire          frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_ready;                             // agent_pipeline_015:in_ready -> frequency_counter_0_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_008_source0_ready;                                                                         // agent_pipeline_016:in_ready -> mux_pipeline_008:out_ready
	wire          agent_pipeline_016_source0_endofpacket;                                                                 // agent_pipeline_016:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_016_source0_valid;                                                                       // agent_pipeline_016:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_016_source0_startofpacket;                                                               // agent_pipeline_016:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] agent_pipeline_016_source0_data;                                                                        // agent_pipeline_016:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] agent_pipeline_016_source0_channel;                                                                     // agent_pipeline_016:out_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_016_source0_ready;                                                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_016:out_ready
	wire          agent_pipeline_017_source0_endofpacket;                                                                 // agent_pipeline_017:out_endofpacket -> id_router_008:sink_endofpacket
	wire          agent_pipeline_017_source0_valid;                                                                       // agent_pipeline_017:out_valid -> id_router_008:sink_valid
	wire          agent_pipeline_017_source0_startofpacket;                                                               // agent_pipeline_017:out_startofpacket -> id_router_008:sink_startofpacket
	wire   [98:0] agent_pipeline_017_source0_data;                                                                        // agent_pipeline_017:out_data -> id_router_008:sink_data
	wire          agent_pipeline_017_source0_ready;                                                                       // id_router_008:sink_ready -> agent_pipeline_017:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_017:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_017:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_017:in_startofpacket
	wire   [98:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_017:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // agent_pipeline_017:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> mux_pipeline:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> mux_pipeline:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> mux_pipeline:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> mux_pipeline:in_data
	wire    [8:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> mux_pipeline:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                                              // mux_pipeline:in_ready -> cmd_xbar_demux:src0_ready
	wire          mux_pipeline_source0_endofpacket;                                                                       // mux_pipeline:out_endofpacket -> agent_pipeline:in_endofpacket
	wire          mux_pipeline_source0_valid;                                                                             // mux_pipeline:out_valid -> agent_pipeline:in_valid
	wire          mux_pipeline_source0_startofpacket;                                                                     // mux_pipeline:out_startofpacket -> agent_pipeline:in_startofpacket
	wire   [98:0] mux_pipeline_source0_data;                                                                              // mux_pipeline:out_data -> agent_pipeline:in_data
	wire    [8:0] mux_pipeline_source0_channel;                                                                           // mux_pipeline:out_channel -> agent_pipeline:in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                        // cmd_xbar_demux:src1_endofpacket -> mux_pipeline_001:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                              // cmd_xbar_demux:src1_valid -> mux_pipeline_001:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                      // cmd_xbar_demux:src1_startofpacket -> mux_pipeline_001:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src1_data;                                                                               // cmd_xbar_demux:src1_data -> mux_pipeline_001:in_data
	wire    [8:0] cmd_xbar_demux_src1_channel;                                                                            // cmd_xbar_demux:src1_channel -> mux_pipeline_001:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                              // mux_pipeline_001:in_ready -> cmd_xbar_demux:src1_ready
	wire          mux_pipeline_001_source0_endofpacket;                                                                   // mux_pipeline_001:out_endofpacket -> agent_pipeline_002:in_endofpacket
	wire          mux_pipeline_001_source0_valid;                                                                         // mux_pipeline_001:out_valid -> agent_pipeline_002:in_valid
	wire          mux_pipeline_001_source0_startofpacket;                                                                 // mux_pipeline_001:out_startofpacket -> agent_pipeline_002:in_startofpacket
	wire   [98:0] mux_pipeline_001_source0_data;                                                                          // mux_pipeline_001:out_data -> agent_pipeline_002:in_data
	wire    [8:0] mux_pipeline_001_source0_channel;                                                                       // mux_pipeline_001:out_channel -> agent_pipeline_002:in_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                        // cmd_xbar_demux:src2_endofpacket -> mux_pipeline_002:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                              // cmd_xbar_demux:src2_valid -> mux_pipeline_002:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                      // cmd_xbar_demux:src2_startofpacket -> mux_pipeline_002:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src2_data;                                                                               // cmd_xbar_demux:src2_data -> mux_pipeline_002:in_data
	wire    [8:0] cmd_xbar_demux_src2_channel;                                                                            // cmd_xbar_demux:src2_channel -> mux_pipeline_002:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                              // mux_pipeline_002:in_ready -> cmd_xbar_demux:src2_ready
	wire          mux_pipeline_002_source0_endofpacket;                                                                   // mux_pipeline_002:out_endofpacket -> width_adapter:in_endofpacket
	wire          mux_pipeline_002_source0_valid;                                                                         // mux_pipeline_002:out_valid -> width_adapter:in_valid
	wire          mux_pipeline_002_source0_startofpacket;                                                                 // mux_pipeline_002:out_startofpacket -> width_adapter:in_startofpacket
	wire   [98:0] mux_pipeline_002_source0_data;                                                                          // mux_pipeline_002:out_data -> width_adapter:in_data
	wire    [8:0] mux_pipeline_002_source0_channel;                                                                       // mux_pipeline_002:out_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                                        // cmd_xbar_demux:src3_endofpacket -> mux_pipeline_003:in_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                              // cmd_xbar_demux:src3_valid -> mux_pipeline_003:in_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                      // cmd_xbar_demux:src3_startofpacket -> mux_pipeline_003:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src3_data;                                                                               // cmd_xbar_demux:src3_data -> mux_pipeline_003:in_data
	wire    [8:0] cmd_xbar_demux_src3_channel;                                                                            // cmd_xbar_demux:src3_channel -> mux_pipeline_003:in_channel
	wire          cmd_xbar_demux_src3_ready;                                                                              // mux_pipeline_003:in_ready -> cmd_xbar_demux:src3_ready
	wire          mux_pipeline_003_source0_endofpacket;                                                                   // mux_pipeline_003:out_endofpacket -> agent_pipeline_006:in_endofpacket
	wire          mux_pipeline_003_source0_valid;                                                                         // mux_pipeline_003:out_valid -> agent_pipeline_006:in_valid
	wire          mux_pipeline_003_source0_startofpacket;                                                                 // mux_pipeline_003:out_startofpacket -> agent_pipeline_006:in_startofpacket
	wire   [98:0] mux_pipeline_003_source0_data;                                                                          // mux_pipeline_003:out_data -> agent_pipeline_006:in_data
	wire    [8:0] mux_pipeline_003_source0_channel;                                                                       // mux_pipeline_003:out_channel -> agent_pipeline_006:in_channel
	wire          cmd_xbar_demux_src4_endofpacket;                                                                        // cmd_xbar_demux:src4_endofpacket -> mux_pipeline_004:in_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                              // cmd_xbar_demux:src4_valid -> mux_pipeline_004:in_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                      // cmd_xbar_demux:src4_startofpacket -> mux_pipeline_004:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src4_data;                                                                               // cmd_xbar_demux:src4_data -> mux_pipeline_004:in_data
	wire    [8:0] cmd_xbar_demux_src4_channel;                                                                            // cmd_xbar_demux:src4_channel -> mux_pipeline_004:in_channel
	wire          cmd_xbar_demux_src4_ready;                                                                              // mux_pipeline_004:in_ready -> cmd_xbar_demux:src4_ready
	wire          mux_pipeline_004_source0_endofpacket;                                                                   // mux_pipeline_004:out_endofpacket -> agent_pipeline_008:in_endofpacket
	wire          mux_pipeline_004_source0_valid;                                                                         // mux_pipeline_004:out_valid -> agent_pipeline_008:in_valid
	wire          mux_pipeline_004_source0_startofpacket;                                                                 // mux_pipeline_004:out_startofpacket -> agent_pipeline_008:in_startofpacket
	wire   [98:0] mux_pipeline_004_source0_data;                                                                          // mux_pipeline_004:out_data -> agent_pipeline_008:in_data
	wire    [8:0] mux_pipeline_004_source0_channel;                                                                       // mux_pipeline_004:out_channel -> agent_pipeline_008:in_channel
	wire          cmd_xbar_demux_src5_endofpacket;                                                                        // cmd_xbar_demux:src5_endofpacket -> mux_pipeline_005:in_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                              // cmd_xbar_demux:src5_valid -> mux_pipeline_005:in_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                      // cmd_xbar_demux:src5_startofpacket -> mux_pipeline_005:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src5_data;                                                                               // cmd_xbar_demux:src5_data -> mux_pipeline_005:in_data
	wire    [8:0] cmd_xbar_demux_src5_channel;                                                                            // cmd_xbar_demux:src5_channel -> mux_pipeline_005:in_channel
	wire          cmd_xbar_demux_src5_ready;                                                                              // mux_pipeline_005:in_ready -> cmd_xbar_demux:src5_ready
	wire          mux_pipeline_005_source0_endofpacket;                                                                   // mux_pipeline_005:out_endofpacket -> width_adapter_002:in_endofpacket
	wire          mux_pipeline_005_source0_valid;                                                                         // mux_pipeline_005:out_valid -> width_adapter_002:in_valid
	wire          mux_pipeline_005_source0_startofpacket;                                                                 // mux_pipeline_005:out_startofpacket -> width_adapter_002:in_startofpacket
	wire   [98:0] mux_pipeline_005_source0_data;                                                                          // mux_pipeline_005:out_data -> width_adapter_002:in_data
	wire    [8:0] mux_pipeline_005_source0_channel;                                                                       // mux_pipeline_005:out_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_src6_endofpacket;                                                                        // cmd_xbar_demux:src6_endofpacket -> mux_pipeline_006:in_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                              // cmd_xbar_demux:src6_valid -> mux_pipeline_006:in_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                      // cmd_xbar_demux:src6_startofpacket -> mux_pipeline_006:in_startofpacket
	wire   [98:0] cmd_xbar_demux_src6_data;                                                                               // cmd_xbar_demux:src6_data -> mux_pipeline_006:in_data
	wire    [8:0] cmd_xbar_demux_src6_channel;                                                                            // cmd_xbar_demux:src6_channel -> mux_pipeline_006:in_channel
	wire          cmd_xbar_demux_src6_ready;                                                                              // mux_pipeline_006:in_ready -> cmd_xbar_demux:src6_ready
	wire          mux_pipeline_006_source0_endofpacket;                                                                   // mux_pipeline_006:out_endofpacket -> agent_pipeline_012:in_endofpacket
	wire          mux_pipeline_006_source0_valid;                                                                         // mux_pipeline_006:out_valid -> agent_pipeline_012:in_valid
	wire          mux_pipeline_006_source0_startofpacket;                                                                 // mux_pipeline_006:out_startofpacket -> agent_pipeline_012:in_startofpacket
	wire   [98:0] mux_pipeline_006_source0_data;                                                                          // mux_pipeline_006:out_data -> agent_pipeline_012:in_data
	wire    [8:0] mux_pipeline_006_source0_channel;                                                                       // mux_pipeline_006:out_channel -> agent_pipeline_012:in_channel
	wire          crosser_out_endofpacket;                                                                                // crosser:out_endofpacket -> mux_pipeline_007:in_endofpacket
	wire          crosser_out_valid;                                                                                      // crosser:out_valid -> mux_pipeline_007:in_valid
	wire          crosser_out_startofpacket;                                                                              // crosser:out_startofpacket -> mux_pipeline_007:in_startofpacket
	wire   [98:0] crosser_out_data;                                                                                       // crosser:out_data -> mux_pipeline_007:in_data
	wire    [8:0] crosser_out_channel;                                                                                    // crosser:out_channel -> mux_pipeline_007:in_channel
	wire          crosser_out_ready;                                                                                      // mux_pipeline_007:in_ready -> crosser:out_ready
	wire          mux_pipeline_007_source0_endofpacket;                                                                   // mux_pipeline_007:out_endofpacket -> agent_pipeline_014:in_endofpacket
	wire          mux_pipeline_007_source0_valid;                                                                         // mux_pipeline_007:out_valid -> agent_pipeline_014:in_valid
	wire          mux_pipeline_007_source0_startofpacket;                                                                 // mux_pipeline_007:out_startofpacket -> agent_pipeline_014:in_startofpacket
	wire   [98:0] mux_pipeline_007_source0_data;                                                                          // mux_pipeline_007:out_data -> agent_pipeline_014:in_data
	wire    [8:0] mux_pipeline_007_source0_channel;                                                                       // mux_pipeline_007:out_channel -> agent_pipeline_014:in_channel
	wire          crosser_001_out_endofpacket;                                                                            // crosser_001:out_endofpacket -> mux_pipeline_008:in_endofpacket
	wire          crosser_001_out_valid;                                                                                  // crosser_001:out_valid -> mux_pipeline_008:in_valid
	wire          crosser_001_out_startofpacket;                                                                          // crosser_001:out_startofpacket -> mux_pipeline_008:in_startofpacket
	wire   [98:0] crosser_001_out_data;                                                                                   // crosser_001:out_data -> mux_pipeline_008:in_data
	wire    [8:0] crosser_001_out_channel;                                                                                // crosser_001:out_channel -> mux_pipeline_008:in_channel
	wire          crosser_001_out_ready;                                                                                  // mux_pipeline_008:in_ready -> crosser_001:out_ready
	wire          mux_pipeline_008_source0_endofpacket;                                                                   // mux_pipeline_008:out_endofpacket -> agent_pipeline_016:in_endofpacket
	wire          mux_pipeline_008_source0_valid;                                                                         // mux_pipeline_008:out_valid -> agent_pipeline_016:in_valid
	wire          mux_pipeline_008_source0_startofpacket;                                                                 // mux_pipeline_008:out_startofpacket -> agent_pipeline_016:in_startofpacket
	wire   [98:0] mux_pipeline_008_source0_data;                                                                          // mux_pipeline_008:out_data -> agent_pipeline_016:in_data
	wire    [8:0] mux_pipeline_008_source0_channel;                                                                       // mux_pipeline_008:out_channel -> agent_pipeline_016:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> mux_pipeline_009:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> mux_pipeline_009:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> mux_pipeline_009:in_startofpacket
	wire   [98:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> mux_pipeline_009:in_data
	wire    [8:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> mux_pipeline_009:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                                              // mux_pipeline_009:in_ready -> rsp_xbar_demux:src0_ready
	wire          mux_pipeline_009_source0_endofpacket;                                                                   // mux_pipeline_009:out_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          mux_pipeline_009_source0_valid;                                                                         // mux_pipeline_009:out_valid -> rsp_xbar_mux:sink0_valid
	wire          mux_pipeline_009_source0_startofpacket;                                                                 // mux_pipeline_009:out_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [98:0] mux_pipeline_009_source0_data;                                                                          // mux_pipeline_009:out_data -> rsp_xbar_mux:sink0_data
	wire    [8:0] mux_pipeline_009_source0_channel;                                                                       // mux_pipeline_009:out_channel -> rsp_xbar_mux:sink0_channel
	wire          mux_pipeline_009_source0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> mux_pipeline_009:out_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> mux_pipeline_010:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> mux_pipeline_010:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> mux_pipeline_010:in_startofpacket
	wire   [98:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> mux_pipeline_010:in_data
	wire    [8:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> mux_pipeline_010:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                          // mux_pipeline_010:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          mux_pipeline_010_source0_endofpacket;                                                                   // mux_pipeline_010:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          mux_pipeline_010_source0_valid;                                                                         // mux_pipeline_010:out_valid -> rsp_xbar_mux:sink1_valid
	wire          mux_pipeline_010_source0_startofpacket;                                                                 // mux_pipeline_010:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [98:0] mux_pipeline_010_source0_data;                                                                          // mux_pipeline_010:out_data -> rsp_xbar_mux:sink1_data
	wire    [8:0] mux_pipeline_010_source0_channel;                                                                       // mux_pipeline_010:out_channel -> rsp_xbar_mux:sink1_channel
	wire          mux_pipeline_010_source0_ready;                                                                         // rsp_xbar_mux:sink1_ready -> mux_pipeline_010:out_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> mux_pipeline_011:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> mux_pipeline_011:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> mux_pipeline_011:in_startofpacket
	wire   [98:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> mux_pipeline_011:in_data
	wire    [8:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> mux_pipeline_011:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                          // mux_pipeline_011:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          mux_pipeline_011_source0_endofpacket;                                                                   // mux_pipeline_011:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          mux_pipeline_011_source0_valid;                                                                         // mux_pipeline_011:out_valid -> rsp_xbar_mux:sink2_valid
	wire          mux_pipeline_011_source0_startofpacket;                                                                 // mux_pipeline_011:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [98:0] mux_pipeline_011_source0_data;                                                                          // mux_pipeline_011:out_data -> rsp_xbar_mux:sink2_data
	wire    [8:0] mux_pipeline_011_source0_channel;                                                                       // mux_pipeline_011:out_channel -> rsp_xbar_mux:sink2_channel
	wire          mux_pipeline_011_source0_ready;                                                                         // rsp_xbar_mux:sink2_ready -> mux_pipeline_011:out_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> mux_pipeline_012:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> mux_pipeline_012:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> mux_pipeline_012:in_startofpacket
	wire   [98:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> mux_pipeline_012:in_data
	wire    [8:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> mux_pipeline_012:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                          // mux_pipeline_012:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          mux_pipeline_012_source0_endofpacket;                                                                   // mux_pipeline_012:out_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          mux_pipeline_012_source0_valid;                                                                         // mux_pipeline_012:out_valid -> rsp_xbar_mux:sink3_valid
	wire          mux_pipeline_012_source0_startofpacket;                                                                 // mux_pipeline_012:out_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire   [98:0] mux_pipeline_012_source0_data;                                                                          // mux_pipeline_012:out_data -> rsp_xbar_mux:sink3_data
	wire    [8:0] mux_pipeline_012_source0_channel;                                                                       // mux_pipeline_012:out_channel -> rsp_xbar_mux:sink3_channel
	wire          mux_pipeline_012_source0_ready;                                                                         // rsp_xbar_mux:sink3_ready -> mux_pipeline_012:out_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> mux_pipeline_013:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> mux_pipeline_013:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> mux_pipeline_013:in_startofpacket
	wire   [98:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> mux_pipeline_013:in_data
	wire    [8:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> mux_pipeline_013:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                          // mux_pipeline_013:in_ready -> rsp_xbar_demux_004:src0_ready
	wire          mux_pipeline_013_source0_endofpacket;                                                                   // mux_pipeline_013:out_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          mux_pipeline_013_source0_valid;                                                                         // mux_pipeline_013:out_valid -> rsp_xbar_mux:sink4_valid
	wire          mux_pipeline_013_source0_startofpacket;                                                                 // mux_pipeline_013:out_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire   [98:0] mux_pipeline_013_source0_data;                                                                          // mux_pipeline_013:out_data -> rsp_xbar_mux:sink4_data
	wire    [8:0] mux_pipeline_013_source0_channel;                                                                       // mux_pipeline_013:out_channel -> rsp_xbar_mux:sink4_channel
	wire          mux_pipeline_013_source0_ready;                                                                         // rsp_xbar_mux:sink4_ready -> mux_pipeline_013:out_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                    // rsp_xbar_demux_005:src0_endofpacket -> mux_pipeline_014:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                          // rsp_xbar_demux_005:src0_valid -> mux_pipeline_014:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                  // rsp_xbar_demux_005:src0_startofpacket -> mux_pipeline_014:in_startofpacket
	wire   [98:0] rsp_xbar_demux_005_src0_data;                                                                           // rsp_xbar_demux_005:src0_data -> mux_pipeline_014:in_data
	wire    [8:0] rsp_xbar_demux_005_src0_channel;                                                                        // rsp_xbar_demux_005:src0_channel -> mux_pipeline_014:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                          // mux_pipeline_014:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          mux_pipeline_014_source0_endofpacket;                                                                   // mux_pipeline_014:out_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          mux_pipeline_014_source0_valid;                                                                         // mux_pipeline_014:out_valid -> rsp_xbar_mux:sink5_valid
	wire          mux_pipeline_014_source0_startofpacket;                                                                 // mux_pipeline_014:out_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire   [98:0] mux_pipeline_014_source0_data;                                                                          // mux_pipeline_014:out_data -> rsp_xbar_mux:sink5_data
	wire    [8:0] mux_pipeline_014_source0_channel;                                                                       // mux_pipeline_014:out_channel -> rsp_xbar_mux:sink5_channel
	wire          mux_pipeline_014_source0_ready;                                                                         // rsp_xbar_mux:sink5_ready -> mux_pipeline_014:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                    // rsp_xbar_demux_006:src0_endofpacket -> mux_pipeline_015:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                          // rsp_xbar_demux_006:src0_valid -> mux_pipeline_015:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                  // rsp_xbar_demux_006:src0_startofpacket -> mux_pipeline_015:in_startofpacket
	wire   [98:0] rsp_xbar_demux_006_src0_data;                                                                           // rsp_xbar_demux_006:src0_data -> mux_pipeline_015:in_data
	wire    [8:0] rsp_xbar_demux_006_src0_channel;                                                                        // rsp_xbar_demux_006:src0_channel -> mux_pipeline_015:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                          // mux_pipeline_015:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          mux_pipeline_015_source0_endofpacket;                                                                   // mux_pipeline_015:out_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          mux_pipeline_015_source0_valid;                                                                         // mux_pipeline_015:out_valid -> rsp_xbar_mux:sink6_valid
	wire          mux_pipeline_015_source0_startofpacket;                                                                 // mux_pipeline_015:out_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire   [98:0] mux_pipeline_015_source0_data;                                                                          // mux_pipeline_015:out_data -> rsp_xbar_mux:sink6_data
	wire    [8:0] mux_pipeline_015_source0_channel;                                                                       // mux_pipeline_015:out_channel -> rsp_xbar_mux:sink6_channel
	wire          mux_pipeline_015_source0_ready;                                                                         // rsp_xbar_mux:sink6_ready -> mux_pipeline_015:out_ready
	wire          crosser_002_out_endofpacket;                                                                            // crosser_002:out_endofpacket -> mux_pipeline_016:in_endofpacket
	wire          crosser_002_out_valid;                                                                                  // crosser_002:out_valid -> mux_pipeline_016:in_valid
	wire          crosser_002_out_startofpacket;                                                                          // crosser_002:out_startofpacket -> mux_pipeline_016:in_startofpacket
	wire   [98:0] crosser_002_out_data;                                                                                   // crosser_002:out_data -> mux_pipeline_016:in_data
	wire    [8:0] crosser_002_out_channel;                                                                                // crosser_002:out_channel -> mux_pipeline_016:in_channel
	wire          crosser_002_out_ready;                                                                                  // mux_pipeline_016:in_ready -> crosser_002:out_ready
	wire          mux_pipeline_016_source0_endofpacket;                                                                   // mux_pipeline_016:out_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          mux_pipeline_016_source0_valid;                                                                         // mux_pipeline_016:out_valid -> rsp_xbar_mux:sink7_valid
	wire          mux_pipeline_016_source0_startofpacket;                                                                 // mux_pipeline_016:out_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire   [98:0] mux_pipeline_016_source0_data;                                                                          // mux_pipeline_016:out_data -> rsp_xbar_mux:sink7_data
	wire    [8:0] mux_pipeline_016_source0_channel;                                                                       // mux_pipeline_016:out_channel -> rsp_xbar_mux:sink7_channel
	wire          mux_pipeline_016_source0_ready;                                                                         // rsp_xbar_mux:sink7_ready -> mux_pipeline_016:out_ready
	wire          crosser_003_out_endofpacket;                                                                            // crosser_003:out_endofpacket -> mux_pipeline_017:in_endofpacket
	wire          crosser_003_out_valid;                                                                                  // crosser_003:out_valid -> mux_pipeline_017:in_valid
	wire          crosser_003_out_startofpacket;                                                                          // crosser_003:out_startofpacket -> mux_pipeline_017:in_startofpacket
	wire   [98:0] crosser_003_out_data;                                                                                   // crosser_003:out_data -> mux_pipeline_017:in_data
	wire    [8:0] crosser_003_out_channel;                                                                                // crosser_003:out_channel -> mux_pipeline_017:in_channel
	wire          crosser_003_out_ready;                                                                                  // mux_pipeline_017:in_ready -> crosser_003:out_ready
	wire          mux_pipeline_017_source0_endofpacket;                                                                   // mux_pipeline_017:out_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          mux_pipeline_017_source0_valid;                                                                         // mux_pipeline_017:out_valid -> rsp_xbar_mux:sink8_valid
	wire          mux_pipeline_017_source0_startofpacket;                                                                 // mux_pipeline_017:out_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire   [98:0] mux_pipeline_017_source0_data;                                                                          // mux_pipeline_017:out_data -> rsp_xbar_mux:sink8_data
	wire    [8:0] mux_pipeline_017_source0_channel;                                                                       // mux_pipeline_017:out_channel -> rsp_xbar_mux:sink8_channel
	wire          mux_pipeline_017_source0_ready;                                                                         // rsp_xbar_mux:sink8_ready -> mux_pipeline_017:out_ready

	mtm_prbs_pattern_generator #(
		.DATA_WIDTH (64),
		.PRBS_WIDTH (32)
	) prbs_pattern_generator (
		.clk            (clk_clk),                                                              //             clock.clk
		.reset          (rst_controller_reset_out_reset),                                       //             reset.reset
		.csr_address    (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_address),    //               csr.address
		.csr_writedata  (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.csr_write      (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_write),      //                  .write
		.csr_readdata   (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.csr_read       (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_read),       //                  .read
		.csr_byteenable (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_byteenable), //                  .byteenable
		.src_data       (prbs_pattern_generator_st_pattern_output_data),                        // st_pattern_output.data
		.src_valid      (prbs_pattern_generator_st_pattern_output_valid),                       //                  .valid
		.src_ready      (prbs_pattern_generator_st_pattern_output_ready)                        //                  .ready
	);

	mtm_prbs_pattern_checker #(
		.DATA_WIDTH (64),
		.PRBS_WIDTH (32)
	) prbs_pattern_checker (
		.clk            (clk_clk),                                                            //            clock.clk
		.reset          (rst_controller_reset_out_reset),                                     //            reset.reset
		.csr_address    (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_address),    //              csr.address
		.csr_writedata  (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_write      (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_readdata   (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.csr_read       (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_byteenable (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_byteenable), //                 .byteenable
		.snk_data       (dma_read_master_data_source_data),                                   // st_pattern_input.data
		.snk_valid      (dma_read_master_data_source_valid),                                  //                 .valid
		.snk_ready      (dma_read_master_data_source_ready)                                   //                 .ready
	);

	write_master #(
		.DATA_WIDTH                     (64),
		.LENGTH_WIDTH                   (31),
		.FIFO_DEPTH                     (128),
		.STRIDE_ENABLE                  (0),
		.BURST_ENABLE                   (1),
		.PACKET_ENABLE                  (0),
		.ERROR_ENABLE                   (0),
		.ERROR_WIDTH                    (8),
		.BYTE_ENABLE_WIDTH              (8),
		.BYTE_ENABLE_WIDTH_LOG2         (3),
		.ADDRESS_WIDTH                  (32),
		.FIFO_DEPTH_LOG2                (7),
		.SYMBOL_WIDTH                   (8),
		.NUMBER_OF_SYMBOLS              (8),
		.NUMBER_OF_SYMBOLS_LOG2         (3),
		.MAX_BURST_COUNT_WIDTH          (6),
		.UNALIGNED_ACCESSES_ENABLE      (0),
		.ONLY_FULL_ACCESS_ENABLE        (1),
		.BURST_WRAPPING_SUPPORT         (0),
		.PROGRAMMABLE_BURST_ENABLE      (0),
		.MAX_BURST_COUNT                (32),
		.FIFO_SPEED_OPTIMIZATION        (1),
		.STRIDE_WIDTH                   (1),
		.ACTUAL_BYTES_TRANSFERRED_WIDTH (32)
	) dma_write_master (
		.clk                (clk_clk),                                     //             Clock.clk
		.reset              (rst_controller_reset_out_reset),              //       Clock_reset.reset
		.master_address     (dma_write_master_address),                    // Data_Write_Master.address
		.master_write       (dma_write_master_write),                      //                  .write
		.master_byteenable  (dma_write_master_byteenable),                 //                  .byteenable
		.master_writedata   (dma_write_master_writedata),                  //                  .writedata
		.master_waitrequest (dma_write_master_waitrequest),                //                  .waitrequest
		.master_burstcount  (dma_write_master_burstcount),                 //                  .burstcount
		.snk_data           (timing_adapter_out_data),                     //         Data_Sink.data
		.snk_valid          (timing_adapter_out_valid),                    //                  .valid
		.snk_ready          (timing_adapter_out_ready),                    //                  .ready
		.snk_command_data   (dispatcher_write_write_command_source_data),  //      Command_Sink.data
		.snk_command_valid  (dispatcher_write_write_command_source_valid), //                  .valid
		.snk_command_ready  (dispatcher_write_write_command_source_ready), //                  .ready
		.src_response_data  (dma_write_master_response_source_data),       //   Response_Source.data
		.src_response_valid (dma_write_master_response_source_valid),      //                  .valid
		.src_response_ready (dma_write_master_response_source_ready),      //                  .ready
		.snk_sop            (1'b0),                                        //       (terminated)
		.snk_eop            (1'b0),                                        //       (terminated)
		.snk_empty          (3'b000),                                      //       (terminated)
		.snk_error          (8'b00000000)                                  //       (terminated)
	);

	dispatcher #(
		.MODE                        (2),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16),
		.CSR_ADDRESS_WIDTH           (3)
	) dispatcher_write (
		.clk                     (clk_clk),                                                                                                                                                                                                                                                               //                clock.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                        //          clock_reset.reset
		.csr_writedata           (dispatcher_write_csr_translator_avalon_anti_slave_0_writedata),                                                                                                                                                                                                         //                  CSR.writedata
		.csr_write               (dispatcher_write_csr_translator_avalon_anti_slave_0_write),                                                                                                                                                                                                             //                     .write
		.csr_byteenable          (dispatcher_write_csr_translator_avalon_anti_slave_0_byteenable),                                                                                                                                                                                                        //                     .byteenable
		.csr_readdata            (dispatcher_write_csr_translator_avalon_anti_slave_0_readdata),                                                                                                                                                                                                          //                     .readdata
		.csr_read                (dispatcher_write_csr_translator_avalon_anti_slave_0_read),                                                                                                                                                                                                              //                     .read
		.csr_address             (dispatcher_write_csr_translator_avalon_anti_slave_0_address),                                                                                                                                                                                                           //                     .address
		.descriptor_write        (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_write),                                                                                                                                                                                                //     Descriptor_Slave.write
		.descriptor_waitrequest  (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_waitrequest),                                                                                                                                                                                          //                     .waitrequest
		.descriptor_writedata    (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_writedata),                                                                                                                                                                                            //                     .writedata
		.descriptor_byteenable   (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_byteenable),                                                                                                                                                                                           //                     .byteenable
		.src_write_master_data   (dispatcher_write_write_command_source_data),                                                                                                                                                                                                                            // Write_Command_Source.data
		.src_write_master_valid  (dispatcher_write_write_command_source_valid),                                                                                                                                                                                                                           //                     .valid
		.src_write_master_ready  (dispatcher_write_write_command_source_ready),                                                                                                                                                                                                                           //                     .ready
		.snk_write_master_data   (dma_write_master_response_source_data),                                                                                                                                                                                                                                 //  Write_Response_Sink.data
		.snk_write_master_valid  (dma_write_master_response_source_valid),                                                                                                                                                                                                                                //                     .valid
		.snk_write_master_ready  (dma_write_master_response_source_ready),                                                                                                                                                                                                                                //                     .ready
		.csr_irq                 (dispatcher_write_csr_irq_irq),                                                                                                                                                                                                                                          //              csr_irq.irq
		.src_response_data       (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_valid      (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_ready      (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_waitrequest (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                                                                                                                                                               //          (terminated)
		.mm_response_address     (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_readdata    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_read        (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.src_read_master_data    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_valid   (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_ready   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_data    (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //          (terminated)
		.snk_read_master_valid   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_ready   ()                                                                                                                                                                                                                                                                       //          (terminated)
	);

	read_master #(
		.DATA_WIDTH                (64),
		.LENGTH_WIDTH              (31),
		.FIFO_DEPTH                (128),
		.STRIDE_ENABLE             (0),
		.BURST_ENABLE              (1),
		.PACKET_ENABLE             (0),
		.ERROR_ENABLE              (0),
		.ERROR_WIDTH               (8),
		.CHANNEL_ENABLE            (0),
		.CHANNEL_WIDTH             (8),
		.BYTE_ENABLE_WIDTH         (8),
		.BYTE_ENABLE_WIDTH_LOG2    (3),
		.ADDRESS_WIDTH             (32),
		.FIFO_DEPTH_LOG2           (7),
		.SYMBOL_WIDTH              (8),
		.NUMBER_OF_SYMBOLS         (8),
		.NUMBER_OF_SYMBOLS_LOG2    (3),
		.MAX_BURST_COUNT_WIDTH     (6),
		.UNALIGNED_ACCESSES_ENABLE (0),
		.ONLY_FULL_ACCESS_ENABLE   (1),
		.BURST_WRAPPING_SUPPORT    (0),
		.PROGRAMMABLE_BURST_ENABLE (0),
		.MAX_BURST_COUNT           (32),
		.FIFO_SPEED_OPTIMIZATION   (1),
		.STRIDE_WIDTH              (1)
	) dma_read_master (
		.clk                  (clk_clk),                                   //            Clock.clk
		.reset                (rst_controller_reset_out_reset),            //      Clock_reset.reset
		.master_address       (dma_read_master_address),                   // Data_Read_Master.address
		.master_read          (dma_read_master_read),                      //                 .read
		.master_byteenable    (dma_read_master_byteenable),                //                 .byteenable
		.master_readdata      (dma_read_master_readdata),                  //                 .readdata
		.master_waitrequest   (dma_read_master_waitrequest),               //                 .waitrequest
		.master_readdatavalid (dma_read_master_readdatavalid),             //                 .readdatavalid
		.master_burstcount    (dma_read_master_burstcount),                //                 .burstcount
		.src_data             (dma_read_master_data_source_data),          //      Data_Source.data
		.src_valid            (dma_read_master_data_source_valid),         //                 .valid
		.src_ready            (dma_read_master_data_source_ready),         //                 .ready
		.snk_command_data     (dispatcher_read_read_command_source_data),  //     Command_Sink.data
		.snk_command_valid    (dispatcher_read_read_command_source_valid), //                 .valid
		.snk_command_ready    (dispatcher_read_read_command_source_ready), //                 .ready
		.src_response_data    (dma_read_master_response_source_data),      //  Response_Source.data
		.src_response_valid   (dma_read_master_response_source_valid),     //                 .valid
		.src_response_ready   (dma_read_master_response_source_ready),     //                 .ready
		.src_sop              (),                                          //      (terminated)
		.src_eop              (),                                          //      (terminated)
		.src_empty            (),                                          //      (terminated)
		.src_error            (),                                          //      (terminated)
		.src_channel          ()                                           //      (terminated)
	);

	dispatcher #(
		.MODE                        (1),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16),
		.CSR_ADDRESS_WIDTH           (3)
	) dispatcher_read (
		.clk                     (clk_clk),                                                                                                                                                                                                                                                               //               clock.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                        //         clock_reset.reset
		.csr_writedata           (dispatcher_read_csr_translator_avalon_anti_slave_0_writedata),                                                                                                                                                                                                          //                 CSR.writedata
		.csr_write               (dispatcher_read_csr_translator_avalon_anti_slave_0_write),                                                                                                                                                                                                              //                    .write
		.csr_byteenable          (dispatcher_read_csr_translator_avalon_anti_slave_0_byteenable),                                                                                                                                                                                                         //                    .byteenable
		.csr_readdata            (dispatcher_read_csr_translator_avalon_anti_slave_0_readdata),                                                                                                                                                                                                           //                    .readdata
		.csr_read                (dispatcher_read_csr_translator_avalon_anti_slave_0_read),                                                                                                                                                                                                               //                    .read
		.csr_address             (dispatcher_read_csr_translator_avalon_anti_slave_0_address),                                                                                                                                                                                                            //                    .address
		.descriptor_write        (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_write),                                                                                                                                                                                                 //    Descriptor_Slave.write
		.descriptor_waitrequest  (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_waitrequest),                                                                                                                                                                                           //                    .waitrequest
		.descriptor_writedata    (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_writedata),                                                                                                                                                                                             //                    .writedata
		.descriptor_byteenable   (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_byteenable),                                                                                                                                                                                            //                    .byteenable
		.src_read_master_data    (dispatcher_read_read_command_source_data),                                                                                                                                                                                                                              // Read_Command_Source.data
		.src_read_master_valid   (dispatcher_read_read_command_source_valid),                                                                                                                                                                                                                             //                    .valid
		.src_read_master_ready   (dispatcher_read_read_command_source_ready),                                                                                                                                                                                                                             //                    .ready
		.snk_read_master_data    (dma_read_master_response_source_data),                                                                                                                                                                                                                                  //  Read_Response_Sink.data
		.snk_read_master_valid   (dma_read_master_response_source_valid),                                                                                                                                                                                                                                 //                    .valid
		.snk_read_master_ready   (dma_read_master_response_source_ready),                                                                                                                                                                                                                                 //                    .ready
		.csr_irq                 (dispatcher_read_csr_irq_irq),                                                                                                                                                                                                                                           //             csr_irq.irq
		.src_response_data       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_response_valid      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_response_ready      (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.mm_response_waitrequest (),                                                                                                                                                                                                                                                                      //         (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                                                                                                                                                               //         (terminated)
		.mm_response_address     (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.mm_response_readdata    (),                                                                                                                                                                                                                                                                      //         (terminated)
		.mm_response_read        (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.src_write_master_data   (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_write_master_valid  (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_write_master_ready  (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.snk_write_master_data   (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.snk_write_master_valid  (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.snk_write_master_ready  ()                                                                                                                                                                                                                                                                       //         (terminated)
	);

	q_sys_mSGDMA_0_timing_adapter timing_adapter (
		.clk       (clk_clk),                                        //   clk.clk
		.reset_n   (~rst_controller_reset_out_reset),                // reset.reset_n
		.in_ready  (prbs_pattern_generator_st_pattern_output_ready), //    in.ready
		.in_valid  (prbs_pattern_generator_st_pattern_output_valid), //      .valid
		.in_data   (prbs_pattern_generator_st_pattern_output_data),  //      .data
		.out_ready (timing_adapter_out_ready),                       //   out.ready
		.out_valid (timing_adapter_out_valid),                       //      .valid
		.out_data  (timing_adapter_out_data)                         //      .data
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (20),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_slv (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mm_bridge_slv_waitrequest),      //    s0.waitrequest
		.s0_readdata      (mm_bridge_slv_readdata),         //      .readdata
		.s0_readdatavalid (mm_bridge_slv_readdatavalid),    //      .readdatavalid
		.s0_burstcount    (mm_bridge_slv_burstcount),       //      .burstcount
		.s0_writedata     (mm_bridge_slv_writedata),        //      .writedata
		.s0_address       (mm_bridge_slv_address),          //      .address
		.s0_write         (mm_bridge_slv_write),            //      .write
		.s0_read          (mm_bridge_slv_read),             //      .read
		.s0_byteenable    (mm_bridge_slv_byteenable),       //      .byteenable
		.s0_debugaccess   (mm_bridge_slv_debugaccess),      //      .debugaccess
		.m0_waitrequest   (mm_bridge_slv_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_slv_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_slv_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_slv_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_slv_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_slv_m0_address),       //      .address
		.m0_write         (mm_bridge_slv_m0_write),         //      .write
		.m0_read          (mm_bridge_slv_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_slv_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_slv_m0_debugaccess)    //      .debugaccess
	);

	status_mon status_mon_0 (
		.slv_read_n        (~status_mon_0_slv_translator_avalon_anti_slave_0_read),       //          slv.read_n
		.slv_write_n       (~status_mon_0_slv_translator_avalon_anti_slave_0_write),      //             .write_n
		.slv_address       (status_mon_0_slv_translator_avalon_anti_slave_0_address),     //             .address
		.slv_cs_n          (~status_mon_0_slv_translator_avalon_anti_slave_0_chipselect), //             .chipselect_n
		.slv_data_write    (status_mon_0_slv_translator_avalon_anti_slave_0_writedata),   //             .writedata
		.slv_data_read     (status_mon_0_slv_translator_avalon_anti_slave_0_readdata),    //             .readdata
		.cal_fail_mon      (status_mon_out_cal_fail_mon),                                 //  conduit_end.export
		.cal_success_mon   (status_mon_out_cal_success_mon),                              //             .export
		.init_done_mon     (status_mon_out_init_done_mon),                                //             .export
		.reset_out_n       (reset_source_reset_n),                                        // reset_source.reset_n
		.slv_clk           (clk_clk),                                                     //        clock.clk
		.slv_reset_n       (~rst_controller_reset_out_reset),                             //      reset_n.reset_n
		.local_init_done   (status_mon_in_local_init_done),                               //       status.local_init_done
		.local_cal_success (status_mon_in_local_cal_success),                             //             .local_cal_success
		.local_cal_fail    (status_mon_in_local_cal_fail)                                 //             .local_cal_fail
	);

	frequency_counter #(
		.SYSTEM_CLK_FREQ_PICO_SEC (20000)
	) frequency_counter_0 (
		.reset_n         (~rst_controller_001_reset_out_reset),                                //          reset.reset_n
		.clk             (clk_0_clk),                                                          //          clock.clk
		.csr_address     (frequency_counter_0_csr_translator_avalon_anti_slave_0_address),     //            csr.address
		.csr_read        (frequency_counter_0_csr_translator_avalon_anti_slave_0_read),        //               .read
		.csr_readdata    (frequency_counter_0_csr_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.csr_waitrequest (frequency_counter_0_csr_translator_avalon_anti_slave_0_waitrequest), //               .waitrequest
		.sample_clk      (clk_clk),                                                            //     sample_clk.clk
		.sample_reset_n  (~rst_controller_002_reset_out_reset)                                 // sample_reset_n.reset_n
	);

	q_sys_mSGDMA_0_timer_0 timer_0 (
		.clk        (clk_0_clk),                                            //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        ()                                                      //   irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (20),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) mm_bridge_slv_m0_translator (
		.clk                   (clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address           (mm_bridge_slv_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (mm_bridge_slv_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (mm_bridge_slv_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (mm_bridge_slv_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (mm_bridge_slv_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (mm_bridge_slv_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (mm_bridge_slv_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (mm_bridge_slv_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (mm_bridge_slv_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (mm_bridge_slv_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (mm_bridge_slv_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (mm_bridge_slv_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (mm_bridge_slv_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (mm_bridge_slv_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (mm_bridge_slv_m0_byteenable),                                         //                          .byteenable
		.av_read               (mm_bridge_slv_m0_read),                                               //                          .read
		.av_readdata           (mm_bridge_slv_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (mm_bridge_slv_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (mm_bridge_slv_m0_write),                                              //                          .write
		.av_writedata          (mm_bridge_slv_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (mm_bridge_slv_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prbs_pattern_generator_csr_translator (
		.clk                   (clk_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prbs_pattern_generator_csr_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dispatcher_write_csr_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dispatcher_write_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dispatcher_write_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dispatcher_write_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dispatcher_write_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dispatcher_write_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (dispatcher_write_csr_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (128),
		.UAV_DATA_W                     (128),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (16),
		.UAV_BYTEENABLE_W               (16),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (5),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (16),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dispatcher_write_descriptor_slave_translator (
		.clk                   (clk_clk),                                                                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                                                        //                    reset.reset
		.uav_address           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address),                                                // avalon_universal_slave_0.address
		.uav_burstcount        (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),                                             //                         .burstcount
		.uav_read              (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read),                                                   //                         .read
		.uav_write             (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write),                                                  //                         .write
		.uav_waitrequest       (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),                                            //                         .waitrequest
		.uav_readdatavalid     (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),                                          //                         .readdatavalid
		.uav_byteenable        (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),                                             //                         .byteenable
		.uav_readdata          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                                               //                         .readdata
		.uav_writedata         (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata),                                              //                         .writedata
		.uav_lock              (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock),                                                   //                         .lock
		.uav_debugaccess       (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),                                            //                         .debugaccess
		.av_write              (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_write),                                                                //      avalon_anti_slave_0.write
		.av_writedata          (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_writedata),                                                            //                         .writedata
		.av_byteenable         (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_byteenable),                                                           //                         .byteenable
		.av_waitrequest        (dispatcher_write_descriptor_slave_translator_avalon_anti_slave_0_waitrequest),                                                          //                         .waitrequest
		.av_address            (),                                                                                                                                      //              (terminated)
		.av_read               (),                                                                                                                                      //              (terminated)
		.av_readdata           (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110101011011101111010101101), //              (terminated)
		.av_begintransfer      (),                                                                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                                                                      //              (terminated)
		.av_lock               (),                                                                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                                                                      //              (terminated)
		.av_clken              (),                                                                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) prbs_pattern_checker_csr_translator (
		.clk                   (clk_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (prbs_pattern_checker_csr_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dispatcher_read_csr_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dispatcher_read_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dispatcher_read_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dispatcher_read_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dispatcher_read_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dispatcher_read_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (dispatcher_read_csr_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (128),
		.UAV_DATA_W                     (128),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (16),
		.UAV_BYTEENABLE_W               (16),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (5),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (16),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dispatcher_read_descriptor_slave_translator (
		.clk                   (clk_clk),                                                                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                                                        //                    reset.reset
		.uav_address           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address),                                                 // avalon_universal_slave_0.address
		.uav_burstcount        (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),                                              //                         .burstcount
		.uav_read              (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read),                                                    //                         .read
		.uav_write             (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write),                                                   //                         .write
		.uav_waitrequest       (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),                                             //                         .waitrequest
		.uav_readdatavalid     (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),                                           //                         .readdatavalid
		.uav_byteenable        (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),                                              //                         .byteenable
		.uav_readdata          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                                                //                         .readdata
		.uav_writedata         (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata),                                               //                         .writedata
		.uav_lock              (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock),                                                    //                         .lock
		.uav_debugaccess       (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),                                             //                         .debugaccess
		.av_write              (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_write),                                                                 //      avalon_anti_slave_0.write
		.av_writedata          (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_writedata),                                                             //                         .writedata
		.av_byteenable         (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_byteenable),                                                            //                         .byteenable
		.av_waitrequest        (dispatcher_read_descriptor_slave_translator_avalon_anti_slave_0_waitrequest),                                                           //                         .waitrequest
		.av_address            (),                                                                                                                                      //              (terminated)
		.av_read               (),                                                                                                                                      //              (terminated)
		.av_readdata           (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110101011011101111010101101), //              (terminated)
		.av_begintransfer      (),                                                                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                                                                      //              (terminated)
		.av_lock               (),                                                                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                                                                      //              (terminated)
		.av_clken              (),                                                                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) status_mon_0_slv_translator (
		.clk                   (clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (status_mon_0_slv_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (status_mon_0_slv_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (status_mon_0_slv_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (status_mon_0_slv_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (status_mon_0_slv_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (status_mon_0_slv_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) frequency_counter_0_csr_translator (
		.clk                   (clk_0_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (frequency_counter_0_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (frequency_counter_0_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (frequency_counter_0_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (frequency_counter_0_csr_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_write              (),                                                                                   //              (terminated)
		.av_writedata          (),                                                                                   //              (terminated)
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_0_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.PKT_BURST_TYPE_H          (76),
		.PKT_BURST_TYPE_L          (75),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_TRANS_EXCLUSIVE       (61),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (78),
		.PKT_DATA_SIDEBAND_L       (78),
		.PKT_QOS_H                 (80),
		.PKT_QOS_L                 (80),
		.PKT_ADDR_SIDEBAND_H       (77),
		.PKT_ADDR_SIDEBAND_L       (77),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (31),
		.CACHE_VALUE               (4'b0000)
	) mm_bridge_slv_m0_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address       (mm_bridge_slv_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (mm_bridge_slv_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (mm_bridge_slv_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (mm_bridge_slv_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (mm_bridge_slv_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (mm_bridge_slv_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (mm_bridge_slv_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (mm_bridge_slv_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (mm_bridge_slv_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (mm_bridge_slv_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (mm_bridge_slv_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                        //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                         //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                      //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                  //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                         //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_source0_ready),                                                                    //              cp.ready
		.cp_valid                (agent_pipeline_source0_valid),                                                                    //                .valid
		.cp_data                 (agent_pipeline_source0_data),                                                                     //                .data
		.cp_startofpacket        (agent_pipeline_source0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (agent_pipeline_source0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (agent_pipeline_source0_channel),                                                                  //                .channel
		.rf_sink_ready           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dispatcher_write_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_002_source0_ready),                                                          //              cp.ready
		.cp_valid                (agent_pipeline_002_source0_valid),                                                          //                .valid
		.cp_data                 (agent_pipeline_002_source0_data),                                                           //                .data
		.cp_startofpacket        (agent_pipeline_002_source0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (agent_pipeline_002_source0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (agent_pipeline_002_source0_channel),                                                        //                .channel
		.rf_sink_ready           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (187),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_ADDR_H                (163),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (164),
		.PKT_TRANS_POSTED          (165),
		.PKT_TRANS_WRITE           (166),
		.PKT_TRANS_READ            (167),
		.PKT_TRANS_LOCK            (168),
		.PKT_SRC_ID_H              (192),
		.PKT_SRC_ID_L              (189),
		.PKT_DEST_ID_H             (196),
		.PKT_DEST_ID_L             (193),
		.PKT_BURSTWRAP_H           (179),
		.PKT_BURSTWRAP_L           (175),
		.PKT_BYTE_CNT_H            (174),
		.PKT_BYTE_CNT_L            (170),
		.PKT_PROTECTION_H          (200),
		.PKT_PROTECTION_L          (198),
		.PKT_RESPONSE_STATUS_H     (206),
		.PKT_RESPONSE_STATUS_L     (205),
		.PKT_BURST_SIZE_H          (182),
		.PKT_BURST_SIZE_L          (180),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (207),
		.AVS_BURSTCOUNT_W          (5),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_004_source0_ready),                                                                       //              cp.ready
		.cp_valid                (agent_pipeline_004_source0_valid),                                                                       //                .valid
		.cp_data                 (agent_pipeline_004_source0_data),                                                                        //                .data
		.cp_startofpacket        (agent_pipeline_004_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (agent_pipeline_004_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (agent_pipeline_004_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (208),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_006_source0_ready),                                                              //              cp.ready
		.cp_valid                (agent_pipeline_006_source0_valid),                                                              //                .valid
		.cp_data                 (agent_pipeline_006_source0_data),                                                               //                .data
		.cp_startofpacket        (agent_pipeline_006_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_006_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (agent_pipeline_006_source0_channel),                                                            //                .channel
		.rf_sink_ready           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dispatcher_read_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_008_source0_ready),                                                         //              cp.ready
		.cp_valid                (agent_pipeline_008_source0_valid),                                                         //                .valid
		.cp_data                 (agent_pipeline_008_source0_data),                                                          //                .data
		.cp_startofpacket        (agent_pipeline_008_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (agent_pipeline_008_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (agent_pipeline_008_source0_channel),                                                       //                .channel
		.rf_sink_ready           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (187),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_ADDR_H                (163),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (164),
		.PKT_TRANS_POSTED          (165),
		.PKT_TRANS_WRITE           (166),
		.PKT_TRANS_READ            (167),
		.PKT_TRANS_LOCK            (168),
		.PKT_SRC_ID_H              (192),
		.PKT_SRC_ID_L              (189),
		.PKT_DEST_ID_H             (196),
		.PKT_DEST_ID_L             (193),
		.PKT_BURSTWRAP_H           (179),
		.PKT_BURSTWRAP_L           (175),
		.PKT_BYTE_CNT_H            (174),
		.PKT_BYTE_CNT_L            (170),
		.PKT_PROTECTION_H          (200),
		.PKT_PROTECTION_L          (198),
		.PKT_RESPONSE_STATUS_H     (206),
		.PKT_RESPONSE_STATUS_L     (205),
		.PKT_BURST_SIZE_H          (182),
		.PKT_BURST_SIZE_L          (180),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (207),
		.AVS_BURSTCOUNT_W          (5),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_010_source0_ready),                                                                      //              cp.ready
		.cp_valid                (agent_pipeline_010_source0_valid),                                                                      //                .valid
		.cp_data                 (agent_pipeline_010_source0_data),                                                                       //                .data
		.cp_startofpacket        (agent_pipeline_010_source0_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (agent_pipeline_010_source0_endofpacket),                                                                //                .endofpacket
		.cp_channel              (agent_pipeline_010_source0_channel),                                                                    //                .channel
		.rf_sink_ready           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (208),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) status_mon_0_slv_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (status_mon_0_slv_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_012_source0_ready),                                                      //              cp.ready
		.cp_valid                (agent_pipeline_012_source0_valid),                                                      //                .valid
		.cp_data                 (agent_pipeline_012_source0_data),                                                       //                .data
		.cp_startofpacket        (agent_pipeline_012_source0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (agent_pipeline_012_source0_endofpacket),                                                //                .endofpacket
		.cp_channel              (agent_pipeline_012_source0_channel),                                                    //                .channel
		.rf_sink_ready           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) frequency_counter_0_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_014_source0_ready),                                                             //              cp.ready
		.cp_valid                (agent_pipeline_014_source0_valid),                                                             //                .valid
		.cp_data                 (agent_pipeline_014_source0_data),                                                              //                .data
		.cp_startofpacket        (agent_pipeline_014_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (agent_pipeline_014_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (agent_pipeline_014_source0_channel),                                                           //                .channel
		.rf_sink_ready           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_0_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_016_source0_ready),                                                //              cp.ready
		.cp_valid                (agent_pipeline_016_source0_valid),                                                //                .valid
		.cp_data                 (agent_pipeline_016_source0_data),                                                 //                .data
		.cp_startofpacket        (agent_pipeline_016_source0_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (agent_pipeline_016_source0_endofpacket),                                          //                .endofpacket
		.cp_channel              (agent_pipeline_016_source0_channel),                                              //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_0_clk),                                                                       //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                        // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	q_sys_mSGDMA_0_addr_router addr_router (
		.sink_ready         (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_bridge_slv_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_src_valid),                                                        //          .valid
		.src_data           (addr_router_src_data),                                                         //          .data
		.src_channel        (addr_router_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                   //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router (
		.sink_ready         (agent_pipeline_001_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_001_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_001_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_001_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_001_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_src_ready),                      //       src.ready
		.src_valid          (id_router_src_valid),                      //          .valid
		.src_data           (id_router_src_data),                       //          .data
		.src_channel        (id_router_src_channel),                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                 //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_001 (
		.sink_ready         (agent_pipeline_003_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_003_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_003_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_003_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_003_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                  //       src.ready
		.src_valid          (id_router_001_src_valid),                  //          .valid
		.src_data           (id_router_001_src_data),                   //          .data
		.src_channel        (id_router_001_src_channel),                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router_002 id_router_002 (
		.sink_ready         (agent_pipeline_005_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_005_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_005_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_005_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_005_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                  //       src.ready
		.src_valid          (id_router_002_src_valid),                  //          .valid
		.src_data           (id_router_002_src_data),                   //          .data
		.src_channel        (id_router_002_src_channel),                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_003 (
		.sink_ready         (agent_pipeline_007_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_007_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_007_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_007_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_007_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                  //       src.ready
		.src_valid          (id_router_003_src_valid),                  //          .valid
		.src_data           (id_router_003_src_data),                   //          .data
		.src_channel        (id_router_003_src_channel),                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_004 (
		.sink_ready         (agent_pipeline_009_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_009_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_009_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_009_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_009_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                  //       src.ready
		.src_valid          (id_router_004_src_valid),                  //          .valid
		.src_data           (id_router_004_src_data),                   //          .data
		.src_channel        (id_router_004_src_channel),                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router_002 id_router_005 (
		.sink_ready         (agent_pipeline_011_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_011_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_011_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_011_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_011_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                  //       src.ready
		.src_valid          (id_router_005_src_valid),                  //          .valid
		.src_data           (id_router_005_src_data),                   //          .data
		.src_channel        (id_router_005_src_channel),                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_006 (
		.sink_ready         (agent_pipeline_013_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_013_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_013_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_013_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_013_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                  //       src.ready
		.src_valid          (id_router_006_src_valid),                  //          .valid
		.src_data           (id_router_006_src_data),                   //          .data
		.src_channel        (id_router_006_src_channel),                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_007 (
		.sink_ready         (agent_pipeline_015_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_015_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_015_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_015_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_015_source0_endofpacket),   //          .endofpacket
		.clk                (clk_0_clk),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                  //       src.ready
		.src_valid          (id_router_007_src_valid),                  //          .valid
		.src_data           (id_router_007_src_data),                   //          .data
		.src_channel        (id_router_007_src_channel),                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)             //          .endofpacket
	);

	q_sys_mSGDMA_0_id_router id_router_008 (
		.sink_ready         (agent_pipeline_017_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_017_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_017_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_017_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_017_source0_endofpacket),   //          .endofpacket
		.clk                (clk_0_clk),                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                  //       src.ready
		.src_valid          (id_router_008_src_valid),                  //          .valid
		.src_data           (id_router_008_src_data),                   //          .data
		.src_channel        (id_router_008_src_channel),                //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)             //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.MAX_OUTSTANDING_RESPONSES (17),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (1),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (62),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                                    //       clk.clk
		.reset                  (rst_controller_reset_out_reset),             // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),                      //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),                      //          .valid
		.cmd_sink_data          (addr_router_src_data),                       //          .data
		.cmd_sink_channel       (addr_router_src_channel),                    //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),              //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),                //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),                      //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),                       //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),                    //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),              //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),                //          .endofpacket
		.cmd_src_valid          (limiter_cmd_src_valid),                      //          .valid
		.rsp_sink_ready         (limiter_pipeline_001_source0_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.rsp_sink_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.rsp_sink_data          (limiter_pipeline_001_source0_data),          //          .data
		.rsp_sink_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),                      //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),                      //          .valid
		.rsp_src_data           (limiter_rsp_src_data),                       //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),                    //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),              //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket)                 //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_0_reset_n),                   // reset_in0.reset
		.clk        (clk_0_clk),                          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_0_reset_n),                   // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_0_clk),                          //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	q_sys_mSGDMA_0_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready         (limiter_pipeline_source0_ready),         //      sink.ready
		.sink_channel       (limiter_pipeline_source0_channel),       //          .channel
		.sink_data          (limiter_pipeline_source0_data),          //          .data
		.sink_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.sink_valid         (limiter_pipeline_source0_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),              //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),               //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),        //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),              //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),              //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),               //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),            //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),        //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),              //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),              //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),               //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),            //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),      //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),        //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),              //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),              //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),               //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),            //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),      //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),        //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),              //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),              //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),               //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),            //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),      //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),        //          .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),              //      src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),              //          .valid
		.src5_data          (cmd_xbar_demux_src5_data),               //          .data
		.src5_channel       (cmd_xbar_demux_src5_channel),            //          .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket),      //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),        //          .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),              //      src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),              //          .valid
		.src6_data          (cmd_xbar_demux_src6_data),               //          .data
		.src6_channel       (cmd_xbar_demux_src6_channel),            //          .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket),      //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket),        //          .endofpacket
		.src7_ready         (cmd_xbar_demux_src7_ready),              //      src7.ready
		.src7_valid         (cmd_xbar_demux_src7_valid),              //          .valid
		.src7_data          (cmd_xbar_demux_src7_data),               //          .data
		.src7_channel       (cmd_xbar_demux_src7_channel),            //          .channel
		.src7_startofpacket (cmd_xbar_demux_src7_startofpacket),      //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_src7_endofpacket),        //          .endofpacket
		.src8_ready         (cmd_xbar_demux_src8_ready),              //      src8.ready
		.src8_valid         (cmd_xbar_demux_src8_valid),              //          .valid
		.src8_data          (cmd_xbar_demux_src8_data),               //          .data
		.src8_channel       (cmd_xbar_demux_src8_channel),            //          .channel
		.src8_startofpacket (cmd_xbar_demux_src8_startofpacket),      //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_src8_endofpacket)         //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_0_clk),                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_0_clk),                             //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	q_sys_mSGDMA_0_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                 //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                 //          .valid
		.src_data            (rsp_xbar_mux_src_data),                  //          .data
		.src_channel         (rsp_xbar_mux_src_channel),               //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),         //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),           //          .endofpacket
		.sink0_ready         (mux_pipeline_009_source0_ready),         //     sink0.ready
		.sink0_valid         (mux_pipeline_009_source0_valid),         //          .valid
		.sink0_channel       (mux_pipeline_009_source0_channel),       //          .channel
		.sink0_data          (mux_pipeline_009_source0_data),          //          .data
		.sink0_startofpacket (mux_pipeline_009_source0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_009_source0_endofpacket),   //          .endofpacket
		.sink1_ready         (mux_pipeline_010_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_010_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_010_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_010_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_010_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_010_source0_endofpacket),   //          .endofpacket
		.sink2_ready         (mux_pipeline_011_source0_ready),         //     sink2.ready
		.sink2_valid         (mux_pipeline_011_source0_valid),         //          .valid
		.sink2_channel       (mux_pipeline_011_source0_channel),       //          .channel
		.sink2_data          (mux_pipeline_011_source0_data),          //          .data
		.sink2_startofpacket (mux_pipeline_011_source0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (mux_pipeline_011_source0_endofpacket),   //          .endofpacket
		.sink3_ready         (mux_pipeline_012_source0_ready),         //     sink3.ready
		.sink3_valid         (mux_pipeline_012_source0_valid),         //          .valid
		.sink3_channel       (mux_pipeline_012_source0_channel),       //          .channel
		.sink3_data          (mux_pipeline_012_source0_data),          //          .data
		.sink3_startofpacket (mux_pipeline_012_source0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (mux_pipeline_012_source0_endofpacket),   //          .endofpacket
		.sink4_ready         (mux_pipeline_013_source0_ready),         //     sink4.ready
		.sink4_valid         (mux_pipeline_013_source0_valid),         //          .valid
		.sink4_channel       (mux_pipeline_013_source0_channel),       //          .channel
		.sink4_data          (mux_pipeline_013_source0_data),          //          .data
		.sink4_startofpacket (mux_pipeline_013_source0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (mux_pipeline_013_source0_endofpacket),   //          .endofpacket
		.sink5_ready         (mux_pipeline_014_source0_ready),         //     sink5.ready
		.sink5_valid         (mux_pipeline_014_source0_valid),         //          .valid
		.sink5_channel       (mux_pipeline_014_source0_channel),       //          .channel
		.sink5_data          (mux_pipeline_014_source0_data),          //          .data
		.sink5_startofpacket (mux_pipeline_014_source0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (mux_pipeline_014_source0_endofpacket),   //          .endofpacket
		.sink6_ready         (mux_pipeline_015_source0_ready),         //     sink6.ready
		.sink6_valid         (mux_pipeline_015_source0_valid),         //          .valid
		.sink6_channel       (mux_pipeline_015_source0_channel),       //          .channel
		.sink6_data          (mux_pipeline_015_source0_data),          //          .data
		.sink6_startofpacket (mux_pipeline_015_source0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (mux_pipeline_015_source0_endofpacket),   //          .endofpacket
		.sink7_ready         (mux_pipeline_016_source0_ready),         //     sink7.ready
		.sink7_valid         (mux_pipeline_016_source0_valid),         //          .valid
		.sink7_channel       (mux_pipeline_016_source0_channel),       //          .channel
		.sink7_data          (mux_pipeline_016_source0_data),          //          .data
		.sink7_startofpacket (mux_pipeline_016_source0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (mux_pipeline_016_source0_endofpacket),   //          .endofpacket
		.sink8_ready         (mux_pipeline_017_source0_ready),         //     sink8.ready
		.sink8_valid         (mux_pipeline_017_source0_valid),         //          .valid
		.sink8_channel       (mux_pipeline_017_source0_channel),       //          .channel
		.sink8_data          (mux_pipeline_017_source0_data),          //          .data
		.sink8_startofpacket (mux_pipeline_017_source0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (mux_pipeline_017_source0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (55),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (66),
		.IN_PKT_BYTE_CNT_L             (62),
		.IN_PKT_TRANS_COMPRESSED_READ  (56),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (67),
		.IN_PKT_BURST_SIZE_H           (74),
		.IN_PKT_BURST_SIZE_L           (72),
		.IN_PKT_RESPONSE_STATUS_H      (98),
		.IN_PKT_RESPONSE_STATUS_L      (97),
		.IN_PKT_TRANS_EXCLUSIVE        (61),
		.IN_PKT_BURST_TYPE_H           (76),
		.IN_PKT_BURST_TYPE_L           (75),
		.IN_ST_DATA_W                  (99),
		.OUT_PKT_ADDR_H                (163),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (174),
		.OUT_PKT_BYTE_CNT_L            (170),
		.OUT_PKT_TRANS_COMPRESSED_READ (164),
		.OUT_PKT_BURST_SIZE_H          (182),
		.OUT_PKT_BURST_SIZE_L          (180),
		.OUT_PKT_RESPONSE_STATUS_H     (206),
		.OUT_PKT_RESPONSE_STATUS_L     (205),
		.OUT_PKT_TRANS_EXCLUSIVE       (169),
		.OUT_PKT_BURST_TYPE_H          (184),
		.OUT_PKT_BURST_TYPE_L          (183),
		.OUT_ST_DATA_W                 (207),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clk_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (mux_pipeline_002_source0_valid),         //      sink.valid
		.in_channel           (mux_pipeline_002_source0_channel),       //          .channel
		.in_startofpacket     (mux_pipeline_002_source0_startofpacket), //          .startofpacket
		.in_endofpacket       (mux_pipeline_002_source0_endofpacket),   //          .endofpacket
		.in_ready             (mux_pipeline_002_source0_ready),         //          .ready
		.in_data              (mux_pipeline_002_source0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),          //       src.endofpacket
		.out_data             (width_adapter_src_data),                 //          .data
		.out_channel          (width_adapter_src_channel),              //          .channel
		.out_valid            (width_adapter_src_valid),                //          .valid
		.out_ready            (width_adapter_src_ready),                //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),        //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (163),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (174),
		.IN_PKT_BYTE_CNT_L             (170),
		.IN_PKT_TRANS_COMPRESSED_READ  (164),
		.IN_PKT_BURSTWRAP_H            (179),
		.IN_PKT_BURSTWRAP_L            (175),
		.IN_PKT_BURST_SIZE_H           (182),
		.IN_PKT_BURST_SIZE_L           (180),
		.IN_PKT_RESPONSE_STATUS_H      (206),
		.IN_PKT_RESPONSE_STATUS_L      (205),
		.IN_PKT_TRANS_EXCLUSIVE        (169),
		.IN_PKT_BURST_TYPE_H           (184),
		.IN_PKT_BURST_TYPE_L           (183),
		.IN_ST_DATA_W                  (207),
		.OUT_PKT_ADDR_H                (55),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (66),
		.OUT_PKT_BYTE_CNT_L            (62),
		.OUT_PKT_TRANS_COMPRESSED_READ (56),
		.OUT_PKT_BURST_SIZE_H          (74),
		.OUT_PKT_BURST_SIZE_L          (72),
		.OUT_PKT_RESPONSE_STATUS_H     (98),
		.OUT_PKT_RESPONSE_STATUS_L     (97),
		.OUT_PKT_TRANS_EXCLUSIVE       (61),
		.OUT_PKT_BURST_TYPE_H          (76),
		.OUT_PKT_BURST_TYPE_L          (75),
		.OUT_ST_DATA_W                 (99),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (55),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (66),
		.IN_PKT_BYTE_CNT_L             (62),
		.IN_PKT_TRANS_COMPRESSED_READ  (56),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (67),
		.IN_PKT_BURST_SIZE_H           (74),
		.IN_PKT_BURST_SIZE_L           (72),
		.IN_PKT_RESPONSE_STATUS_H      (98),
		.IN_PKT_RESPONSE_STATUS_L      (97),
		.IN_PKT_TRANS_EXCLUSIVE        (61),
		.IN_PKT_BURST_TYPE_H           (76),
		.IN_PKT_BURST_TYPE_L           (75),
		.IN_ST_DATA_W                  (99),
		.OUT_PKT_ADDR_H                (163),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (174),
		.OUT_PKT_BYTE_CNT_L            (170),
		.OUT_PKT_TRANS_COMPRESSED_READ (164),
		.OUT_PKT_BURST_SIZE_H          (182),
		.OUT_PKT_BURST_SIZE_L          (180),
		.OUT_PKT_RESPONSE_STATUS_H     (206),
		.OUT_PKT_RESPONSE_STATUS_L     (205),
		.OUT_PKT_TRANS_EXCLUSIVE       (169),
		.OUT_PKT_BURST_TYPE_H          (184),
		.OUT_PKT_BURST_TYPE_L          (183),
		.OUT_ST_DATA_W                 (207),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (clk_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (mux_pipeline_005_source0_valid),         //      sink.valid
		.in_channel           (mux_pipeline_005_source0_channel),       //          .channel
		.in_startofpacket     (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.in_endofpacket       (mux_pipeline_005_source0_endofpacket),   //          .endofpacket
		.in_ready             (mux_pipeline_005_source0_ready),         //          .ready
		.in_data              (mux_pipeline_005_source0_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_002_src_data),             //          .data
		.out_channel          (width_adapter_002_src_channel),          //          .channel
		.out_valid            (width_adapter_002_src_valid),            //          .valid
		.out_ready            (width_adapter_002_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (163),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (174),
		.IN_PKT_BYTE_CNT_L             (170),
		.IN_PKT_TRANS_COMPRESSED_READ  (164),
		.IN_PKT_BURSTWRAP_H            (179),
		.IN_PKT_BURSTWRAP_L            (175),
		.IN_PKT_BURST_SIZE_H           (182),
		.IN_PKT_BURST_SIZE_L           (180),
		.IN_PKT_RESPONSE_STATUS_H      (206),
		.IN_PKT_RESPONSE_STATUS_L      (205),
		.IN_PKT_TRANS_EXCLUSIVE        (169),
		.IN_PKT_BURST_TYPE_H           (184),
		.IN_PKT_BURST_TYPE_L           (183),
		.IN_ST_DATA_W                  (207),
		.OUT_PKT_ADDR_H                (55),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (66),
		.OUT_PKT_BYTE_CNT_L            (62),
		.OUT_PKT_TRANS_COMPRESSED_READ (56),
		.OUT_PKT_BURST_SIZE_H          (74),
		.OUT_PKT_BURST_SIZE_L          (72),
		.OUT_PKT_RESPONSE_STATUS_H     (98),
		.OUT_PKT_RESPONSE_STATUS_L     (97),
		.OUT_PKT_TRANS_EXCLUSIVE       (61),
		.OUT_PKT_BURST_TYPE_H          (76),
		.OUT_PKT_BURST_TYPE_L          (75),
		.OUT_ST_DATA_W                 (99),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_005_src_valid),             //      sink.valid
		.in_channel           (id_router_005_src_channel),           //          .channel
		.in_startofpacket     (id_router_005_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_005_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_005_src_ready),             //          .ready
		.in_data              (id_router_005_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_0_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src7_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src7_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src7_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src7_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_0_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src8_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src8_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src8_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src8_data),           //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk_0_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_0_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (limiter_cmd_src_ready),                  //     sink0.ready
		.in_valid          (limiter_cmd_src_valid),                  //          .valid
		.in_startofpacket  (limiter_cmd_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (limiter_cmd_src_endofpacket),            //          .endofpacket
		.in_data           (limiter_cmd_src_data),                   //          .data
		.in_channel        (limiter_cmd_src_channel),                //          .channel
		.out_ready         (limiter_pipeline_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_source0_data),          //          .data
		.out_channel       (limiter_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_001 (
		.clk               (clk_clk),                                    //       cr0.clk
		.reset             (rst_controller_reset_out_reset),             // cr0_reset.reset
		.in_ready          (rsp_xbar_mux_src_ready),                     //     sink0.ready
		.in_valid          (rsp_xbar_mux_src_valid),                     //          .valid
		.in_startofpacket  (rsp_xbar_mux_src_startofpacket),             //          .startofpacket
		.in_endofpacket    (rsp_xbar_mux_src_endofpacket),               //          .endofpacket
		.in_data           (rsp_xbar_mux_src_data),                      //          .data
		.in_channel        (rsp_xbar_mux_src_channel),                   //          .channel
		.out_ready         (limiter_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_001_source0_data),          //          .data
		.out_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline (
		.clk               (clk_clk),                              //       cr0.clk
		.reset             (rst_controller_reset_out_reset),       // cr0_reset.reset
		.in_ready          (mux_pipeline_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_source0_data),            //          .data
		.in_channel        (mux_pipeline_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_source0_data),          //          .data
		.out_channel       (agent_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.out_error         (),                                     // (terminated)
		.in_error          (1'b0)                                  // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_001 (
		.clk               (clk_clk),                                                                               //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                        // cr0_reset.reset
		.in_ready          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (prbs_pattern_generator_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_001_source0_ready),                                                      //   source0.ready
		.out_valid         (agent_pipeline_001_source0_valid),                                                      //          .valid
		.out_startofpacket (agent_pipeline_001_source0_startofpacket),                                              //          .startofpacket
		.out_endofpacket   (agent_pipeline_001_source0_endofpacket),                                                //          .endofpacket
		.out_data          (agent_pipeline_001_source0_data),                                                       //          .data
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_channel       (),                                                                                      // (terminated)
		.in_channel        (1'b0)                                                                                   // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_002 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (mux_pipeline_001_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_001_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_001_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_001_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_001_source0_data),            //          .data
		.in_channel        (mux_pipeline_001_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_002_source0_data),          //          .data
		.out_channel       (agent_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_003 (
		.clk               (clk_clk),                                                                         //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                  // cr0_reset.reset
		.in_ready          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (dispatcher_write_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_003_source0_ready),                                                //   source0.ready
		.out_valid         (agent_pipeline_003_source0_valid),                                                //          .valid
		.out_startofpacket (agent_pipeline_003_source0_startofpacket),                                        //          .startofpacket
		.out_endofpacket   (agent_pipeline_003_source0_endofpacket),                                          //          .endofpacket
		.out_data          (agent_pipeline_003_source0_data),                                                 //          .data
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_channel       (),                                                                                // (terminated)
		.in_channel        (1'b0)                                                                             // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (207),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_004 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (width_adapter_src_ready),                  //     sink0.ready
		.in_valid          (width_adapter_src_valid),                  //          .valid
		.in_startofpacket  (width_adapter_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (width_adapter_src_endofpacket),            //          .endofpacket
		.in_data           (width_adapter_src_data),                   //          .data
		.in_channel        (width_adapter_src_channel),                //          .channel
		.out_ready         (agent_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_004_source0_data),          //          .data
		.out_channel       (agent_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (207),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_005 (
		.clk               (clk_clk),                                                                                      //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                               // cr0_reset.reset
		.in_ready          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (dispatcher_write_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_005_source0_ready),                                                             //   source0.ready
		.out_valid         (agent_pipeline_005_source0_valid),                                                             //          .valid
		.out_startofpacket (agent_pipeline_005_source0_startofpacket),                                                     //          .startofpacket
		.out_endofpacket   (agent_pipeline_005_source0_endofpacket),                                                       //          .endofpacket
		.out_data          (agent_pipeline_005_source0_data),                                                              //          .data
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_channel       (),                                                                                             // (terminated)
		.in_channel        (1'b0)                                                                                          // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_006 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (mux_pipeline_003_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_003_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_003_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_003_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_003_source0_data),            //          .data
		.in_channel        (mux_pipeline_003_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_006_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_006_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_006_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_006_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_006_source0_data),          //          .data
		.out_channel       (agent_pipeline_006_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_007 (
		.clk               (clk_clk),                                                                             //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                      // cr0_reset.reset
		.in_ready          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (prbs_pattern_checker_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_007_source0_ready),                                                    //   source0.ready
		.out_valid         (agent_pipeline_007_source0_valid),                                                    //          .valid
		.out_startofpacket (agent_pipeline_007_source0_startofpacket),                                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_007_source0_endofpacket),                                              //          .endofpacket
		.out_data          (agent_pipeline_007_source0_data),                                                     //          .data
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_channel       (),                                                                                    // (terminated)
		.in_channel        (1'b0)                                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_008 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (mux_pipeline_004_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_004_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_004_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_004_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_004_source0_data),            //          .data
		.in_channel        (mux_pipeline_004_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_008_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_008_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_008_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_008_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_008_source0_data),          //          .data
		.out_channel       (agent_pipeline_008_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_009 (
		.clk               (clk_clk),                                                                        //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                 // cr0_reset.reset
		.in_ready          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (dispatcher_read_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_009_source0_ready),                                               //   source0.ready
		.out_valid         (agent_pipeline_009_source0_valid),                                               //          .valid
		.out_startofpacket (agent_pipeline_009_source0_startofpacket),                                       //          .startofpacket
		.out_endofpacket   (agent_pipeline_009_source0_endofpacket),                                         //          .endofpacket
		.out_data          (agent_pipeline_009_source0_data),                                                //          .data
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_channel       (),                                                                               // (terminated)
		.in_channel        (1'b0)                                                                            // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (207),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_010 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (width_adapter_002_src_ready),              //     sink0.ready
		.in_valid          (width_adapter_002_src_valid),              //          .valid
		.in_startofpacket  (width_adapter_002_src_startofpacket),      //          .startofpacket
		.in_endofpacket    (width_adapter_002_src_endofpacket),        //          .endofpacket
		.in_data           (width_adapter_002_src_data),               //          .data
		.in_channel        (width_adapter_002_src_channel),            //          .channel
		.out_ready         (agent_pipeline_010_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_010_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_010_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_010_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_010_source0_data),          //          .data
		.out_channel       (agent_pipeline_010_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (207),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_011 (
		.clk               (clk_clk),                                                                                     //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                              // cr0_reset.reset
		.in_ready          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (dispatcher_read_descriptor_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_011_source0_ready),                                                            //   source0.ready
		.out_valid         (agent_pipeline_011_source0_valid),                                                            //          .valid
		.out_startofpacket (agent_pipeline_011_source0_startofpacket),                                                    //          .startofpacket
		.out_endofpacket   (agent_pipeline_011_source0_endofpacket),                                                      //          .endofpacket
		.out_data          (agent_pipeline_011_source0_data),                                                             //          .data
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_channel       (),                                                                                            // (terminated)
		.in_channel        (1'b0)                                                                                         // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_012 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (mux_pipeline_006_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_006_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_006_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_006_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_006_source0_data),            //          .data
		.in_channel        (mux_pipeline_006_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_012_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_012_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_012_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_012_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_012_source0_data),          //          .data
		.out_channel       (agent_pipeline_012_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_013 (
		.clk               (clk_clk),                                                                     //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                              // cr0_reset.reset
		.in_ready          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (status_mon_0_slv_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_013_source0_ready),                                            //   source0.ready
		.out_valid         (agent_pipeline_013_source0_valid),                                            //          .valid
		.out_startofpacket (agent_pipeline_013_source0_startofpacket),                                    //          .startofpacket
		.out_endofpacket   (agent_pipeline_013_source0_endofpacket),                                      //          .endofpacket
		.out_data          (agent_pipeline_013_source0_data),                                             //          .data
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_channel       (),                                                                            // (terminated)
		.in_channel        (1'b0)                                                                         // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_014 (
		.clk               (clk_0_clk),                                //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),       // cr0_reset.reset
		.in_ready          (mux_pipeline_007_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_007_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_007_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_007_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_007_source0_data),            //          .data
		.in_channel        (mux_pipeline_007_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_014_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_014_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_014_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_014_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_014_source0_data),          //          .data
		.out_channel       (agent_pipeline_014_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_015 (
		.clk               (clk_0_clk),                                                                          //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // cr0_reset.reset
		.in_ready          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (frequency_counter_0_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_015_source0_ready),                                                   //   source0.ready
		.out_valid         (agent_pipeline_015_source0_valid),                                                   //          .valid
		.out_startofpacket (agent_pipeline_015_source0_startofpacket),                                           //          .startofpacket
		.out_endofpacket   (agent_pipeline_015_source0_endofpacket),                                             //          .endofpacket
		.out_data          (agent_pipeline_015_source0_data),                                                    //          .data
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_channel       (),                                                                                   // (terminated)
		.in_channel        (1'b0)                                                                                // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_016 (
		.clk               (clk_0_clk),                                //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),       // cr0_reset.reset
		.in_ready          (mux_pipeline_008_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_008_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_008_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_008_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_008_source0_data),            //          .data
		.in_channel        (mux_pipeline_008_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_016_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_016_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_016_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_016_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_016_source0_data),          //          .data
		.out_channel       (agent_pipeline_016_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_017 (
		.clk               (clk_0_clk),                                                             //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),                                    // cr0_reset.reset
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_017_source0_ready),                                      //   source0.ready
		.out_valid         (agent_pipeline_017_source0_valid),                                      //          .valid
		.out_startofpacket (agent_pipeline_017_source0_startofpacket),                              //          .startofpacket
		.out_endofpacket   (agent_pipeline_017_source0_endofpacket),                                //          .endofpacket
		.out_data          (agent_pipeline_017_source0_data),                                       //          .data
		.in_empty          (1'b0),                                                                  // (terminated)
		.out_empty         (),                                                                      // (terminated)
		.out_error         (),                                                                      // (terminated)
		.in_error          (1'b0),                                                                  // (terminated)
		.out_channel       (),                                                                      // (terminated)
		.in_channel        (1'b0)                                                                   // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline (
		.clk               (clk_clk),                            //       cr0.clk
		.reset             (rst_controller_reset_out_reset),     // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_src0_data),           //          .data
		.in_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_source0_data),          //          .data
		.out_channel       (mux_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                               // (terminated)
		.out_empty         (),                                   // (terminated)
		.out_error         (),                                   // (terminated)
		.in_error          (1'b0)                                // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_001 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src1_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src1_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src1_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src1_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src1_data),               //          .data
		.in_channel        (cmd_xbar_demux_src1_channel),            //          .channel
		.out_ready         (mux_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_001_source0_data),          //          .data
		.out_channel       (mux_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_002 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src2_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src2_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src2_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src2_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src2_data),               //          .data
		.in_channel        (cmd_xbar_demux_src2_channel),            //          .channel
		.out_ready         (mux_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_002_source0_data),          //          .data
		.out_channel       (mux_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_003 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src3_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src3_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src3_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src3_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src3_data),               //          .data
		.in_channel        (cmd_xbar_demux_src3_channel),            //          .channel
		.out_ready         (mux_pipeline_003_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_003_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_003_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_003_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_003_source0_data),          //          .data
		.out_channel       (mux_pipeline_003_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_004 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src4_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src4_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src4_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src4_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src4_data),               //          .data
		.in_channel        (cmd_xbar_demux_src4_channel),            //          .channel
		.out_ready         (mux_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_004_source0_data),          //          .data
		.out_channel       (mux_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_005 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src5_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src5_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src5_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src5_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src5_data),               //          .data
		.in_channel        (cmd_xbar_demux_src5_channel),            //          .channel
		.out_ready         (mux_pipeline_005_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_005_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_005_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_005_source0_data),          //          .data
		.out_channel       (mux_pipeline_005_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_006 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src6_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src6_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src6_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src6_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src6_data),               //          .data
		.in_channel        (cmd_xbar_demux_src6_channel),            //          .channel
		.out_ready         (mux_pipeline_006_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_006_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_006_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_006_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_006_source0_data),          //          .data
		.out_channel       (mux_pipeline_006_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_007 (
		.clk               (clk_0_clk),                              //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_out_ready),                      //     sink0.ready
		.in_valid          (crosser_out_valid),                      //          .valid
		.in_startofpacket  (crosser_out_startofpacket),              //          .startofpacket
		.in_endofpacket    (crosser_out_endofpacket),                //          .endofpacket
		.in_data           (crosser_out_data),                       //          .data
		.in_channel        (crosser_out_channel),                    //          .channel
		.out_ready         (mux_pipeline_007_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_007_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_007_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_007_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_007_source0_data),          //          .data
		.out_channel       (mux_pipeline_007_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_008 (
		.clk               (clk_0_clk),                              //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_001_out_ready),                  //     sink0.ready
		.in_valid          (crosser_001_out_valid),                  //          .valid
		.in_startofpacket  (crosser_001_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_001_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_001_out_data),                   //          .data
		.in_channel        (crosser_001_out_channel),                //          .channel
		.out_ready         (mux_pipeline_008_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_008_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_008_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_008_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_008_source0_data),          //          .data
		.out_channel       (mux_pipeline_008_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_009 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),              //     sink0.ready
		.in_valid          (rsp_xbar_demux_src0_valid),              //          .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),        //          .endofpacket
		.in_data           (rsp_xbar_demux_src0_data),               //          .data
		.in_channel        (rsp_xbar_demux_src0_channel),            //          .channel
		.out_ready         (mux_pipeline_009_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_009_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_009_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_009_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_009_source0_data),          //          .data
		.out_channel       (mux_pipeline_009_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_010 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_001_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_001_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_001_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_001_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_010_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_010_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_010_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_010_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_010_source0_data),          //          .data
		.out_channel       (mux_pipeline_010_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_011 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_002_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_002_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_002_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_002_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_011_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_011_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_011_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_011_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_011_source0_data),          //          .data
		.out_channel       (mux_pipeline_011_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_012 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_003_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_003_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_003_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_003_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_012_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_012_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_012_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_012_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_012_source0_data),          //          .data
		.out_channel       (mux_pipeline_012_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_013 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_004_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_004_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_013_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_013_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_013_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_013_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_013_source0_data),          //          .data
		.out_channel       (mux_pipeline_013_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_014 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_005_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_005_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_005_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_005_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_005_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_014_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_014_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_014_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_014_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_014_source0_data),          //          .data
		.out_channel       (mux_pipeline_014_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_015 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_006_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_006_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_015_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_015_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_015_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_015_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_015_source0_data),          //          .data
		.out_channel       (mux_pipeline_015_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_016 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (crosser_002_out_ready),                  //     sink0.ready
		.in_valid          (crosser_002_out_valid),                  //          .valid
		.in_startofpacket  (crosser_002_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_002_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_002_out_data),                   //          .data
		.in_channel        (crosser_002_out_channel),                //          .channel
		.out_ready         (mux_pipeline_016_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_016_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_016_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_016_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_016_source0_data),          //          .data
		.out_channel       (mux_pipeline_016_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (99),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (9),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_017 (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),         // cr0_reset.reset
		.in_ready          (crosser_003_out_ready),                  //     sink0.ready
		.in_valid          (crosser_003_out_valid),                  //          .valid
		.in_startofpacket  (crosser_003_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_003_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_003_out_data),                   //          .data
		.in_channel        (crosser_003_out_channel),                //          .channel
		.out_ready         (mux_pipeline_017_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_017_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_017_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_017_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_017_source0_data),          //          .data
		.out_channel       (mux_pipeline_017_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

endmodule
