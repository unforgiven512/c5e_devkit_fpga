// q_sys.v

// Generated using ACDS version 12.1sp1 243 at 2013.02.13.11:10:28

`timescale 1 ps / 1 ps
module q_sys (
		input  wire        oct_rzqin,                                     //                                oct.rzqin
		input  wire        reset_50_reset_n,                              //                           reset_50.reset_n
		output wire        msgdma_0_status_mon_out_cal_fail_mon,          //            msgdma_0_status_mon_out.cal_fail_mon
		output wire        msgdma_0_status_mon_out_cal_success_mon,       //                                   .cal_success_mon
		output wire        msgdma_0_status_mon_out_init_done_mon,         //                                   .init_done_mon
		input  wire        reset_reset_n,                                 //                              reset.reset_n
		input  wire        clk_50_clk,                                    //                             clk_50.clk
		input  wire        clk_clk,                                       //                                clk.clk
		output wire        master_driver_msgdma_0_conduit_end_error_mon,  // master_driver_msgdma_0_conduit_end.error_mon
		output wire        master_driver_msgdma_0_conduit_end_status_mon, //                                   .status_mon
		output wire [9:0]  memory_mem_ca,                                 //                             memory.mem_ca
		output wire [0:0]  memory_mem_ck,                                 //                                   .mem_ck
		output wire [0:0]  memory_mem_ck_n,                               //                                   .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                //                                   .mem_cke
		output wire [0:0]  memory_mem_cs_n,                               //                                   .mem_cs_n
		output wire [1:0]  memory_mem_dm,                                 //                                   .mem_dm
		inout  wire [15:0] memory_mem_dq,                                 //                                   .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                                //                                   .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n                               //                                   .mem_dqs_n
	);

	wire          mem_if_lpddr2_emif_0_afi_clk_clk;                                                                   // mem_if_lpddr2_emif_0:afi_clk -> [addr_router_002:clk, addr_router_003:clk, agent_pipeline_004:clk, agent_pipeline_005:clk, agent_pipeline_006:clk, agent_pipeline_007:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, crosser:out_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, id_router_002:clk, id_router_003:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mSGDMA_0:clk_clk, mSGDMA_0_dma_read_master_translator:clk, mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:clk, mSGDMA_0_dma_write_master_translator:clk, mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:clk, mSGDMA_0_mm_bridge_slv_translator:clk, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:clk, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, mem_if_lpddr2_emif_0_avl_translator:clk, mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:clk, mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, mux_pipeline_002:clk, mux_pipeline_003:clk, mux_pipeline_008:clk, mux_pipeline_009:clk, mux_pipeline_010:clk, mux_pipeline_011:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rst_controller_005:clk, rst_controller_006:clk]
	wire          mem_if_lpddr2_emif_0_status_local_cal_fail;                                                         // mem_if_lpddr2_emif_0:local_cal_fail -> mSGDMA_0:status_mon_in_local_cal_fail
	wire          mem_if_lpddr2_emif_0_status_local_cal_success;                                                      // mem_if_lpddr2_emif_0:local_cal_success -> mSGDMA_0:status_mon_in_local_cal_success
	wire          mem_if_lpddr2_emif_0_status_local_init_done;                                                        // mem_if_lpddr2_emif_0:local_init_done -> mSGDMA_0:status_mon_in_local_init_done
	wire          master_0_master_waitrequest;                                                                        // master_0_master_translator:av_waitrequest -> master_0:master_waitrequest
	wire   [31:0] master_0_master_writedata;                                                                          // master_0:master_writedata -> master_0_master_translator:av_writedata
	wire   [31:0] master_0_master_address;                                                                            // master_0:master_address -> master_0_master_translator:av_address
	wire          master_0_master_write;                                                                              // master_0:master_write -> master_0_master_translator:av_write
	wire          master_0_master_read;                                                                               // master_0:master_read -> master_0_master_translator:av_read
	wire   [31:0] master_0_master_readdata;                                                                           // master_0_master_translator:av_readdata -> master_0:master_readdata
	wire    [3:0] master_0_master_byteenable;                                                                         // master_0:master_byteenable -> master_0_master_translator:av_byteenable
	wire          master_0_master_readdatavalid;                                                                      // master_0_master_translator:av_readdatavalid -> master_0:master_readdatavalid
	wire          master_driver_msgdma_0_avalon_master_waitrequest;                                                   // master_driver_msgdma_0_avalon_master_translator:av_waitrequest -> master_driver_msgdma_0:waitrequest_in
	wire   [31:0] master_driver_msgdma_0_avalon_master_writedata;                                                     // master_driver_msgdma_0:data_write -> master_driver_msgdma_0_avalon_master_translator:av_writedata
	wire   [31:0] master_driver_msgdma_0_avalon_master_address;                                                       // master_driver_msgdma_0:address -> master_driver_msgdma_0_avalon_master_translator:av_address
	wire          master_driver_msgdma_0_avalon_master_chipselect;                                                    // master_driver_msgdma_0:csn -> master_driver_msgdma_0_avalon_master_translator:av_chipselect
	wire          master_driver_msgdma_0_avalon_master_write;                                                         // master_driver_msgdma_0:wen -> master_driver_msgdma_0_avalon_master_translator:av_write
	wire          master_driver_msgdma_0_avalon_master_read;                                                          // master_driver_msgdma_0:oen -> master_driver_msgdma_0_avalon_master_translator:av_read
	wire   [31:0] master_driver_msgdma_0_avalon_master_readdata;                                                      // master_driver_msgdma_0_avalon_master_translator:av_readdata -> master_driver_msgdma_0:data_read
	wire    [3:0] master_driver_msgdma_0_avalon_master_byteenable;                                                    // master_driver_msgdma_0:be -> master_driver_msgdma_0_avalon_master_translator:av_byteenable
	wire          master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_waitrequest;                              // master_driver_msgdma_0:csr_waitrequest -> master_driver_msgdma_0_csr_translator:av_waitrequest
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_writedata;                                // master_driver_msgdma_0_csr_translator:av_writedata -> master_driver_msgdma_0:csr_writedata
	wire    [3:0] master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_address;                                  // master_driver_msgdma_0_csr_translator:av_address -> master_driver_msgdma_0:csr_address
	wire          master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_write;                                    // master_driver_msgdma_0_csr_translator:av_write -> master_driver_msgdma_0:csr_write
	wire          master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_read;                                     // master_driver_msgdma_0_csr_translator:av_read -> master_driver_msgdma_0:csr_read
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_readdata;                                 // master_driver_msgdma_0:csr_readdata -> master_driver_msgdma_0_csr_translator:av_readdata
	wire    [1:0] product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // product_info_0_avalon_slave_0_translator:av_address -> product_info_0:av_address
	wire          product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                            // product_info_0_avalon_slave_0_translator:av_chipselect -> product_info_0:chipselect_n
	wire          product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                  // product_info_0_avalon_slave_0_translator:av_read -> product_info_0:read_n
	wire   [31:0] product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // product_info_0:av_data_read -> product_info_0_avalon_slave_0_translator:av_readdata
	wire          msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_waitrequest;                                  // mSGDMA_0:mm_bridge_slv_waitrequest -> mSGDMA_0_mm_bridge_slv_translator:av_waitrequest
	wire    [0:0] msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_burstcount;                                   // mSGDMA_0_mm_bridge_slv_translator:av_burstcount -> mSGDMA_0:mm_bridge_slv_burstcount
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_writedata;                                    // mSGDMA_0_mm_bridge_slv_translator:av_writedata -> mSGDMA_0:mm_bridge_slv_writedata
	wire   [19:0] msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_address;                                      // mSGDMA_0_mm_bridge_slv_translator:av_address -> mSGDMA_0:mm_bridge_slv_address
	wire          msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_write;                                        // mSGDMA_0_mm_bridge_slv_translator:av_write -> mSGDMA_0:mm_bridge_slv_write
	wire          msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_read;                                         // mSGDMA_0_mm_bridge_slv_translator:av_read -> mSGDMA_0:mm_bridge_slv_read
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdata;                                     // mSGDMA_0:mm_bridge_slv_readdata -> mSGDMA_0_mm_bridge_slv_translator:av_readdata
	wire          msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_debugaccess;                                  // mSGDMA_0_mm_bridge_slv_translator:av_debugaccess -> mSGDMA_0:mm_bridge_slv_debugaccess
	wire          msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdatavalid;                                // mSGDMA_0:mm_bridge_slv_readdatavalid -> mSGDMA_0_mm_bridge_slv_translator:av_readdatavalid
	wire    [3:0] msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_byteenable;                                   // mSGDMA_0_mm_bridge_slv_translator:av_byteenable -> mSGDMA_0:mm_bridge_slv_byteenable
	wire    [5:0] msgdma_0_dma_read_master_burstcount;                                                                // mSGDMA_0:dma_read_master_burstcount -> mSGDMA_0_dma_read_master_translator:av_burstcount
	wire          msgdma_0_dma_read_master_waitrequest;                                                               // mSGDMA_0_dma_read_master_translator:av_waitrequest -> mSGDMA_0:dma_read_master_waitrequest
	wire   [31:0] msgdma_0_dma_read_master_address;                                                                   // mSGDMA_0:dma_read_master_address -> mSGDMA_0_dma_read_master_translator:av_address
	wire          msgdma_0_dma_read_master_read;                                                                      // mSGDMA_0:dma_read_master_read -> mSGDMA_0_dma_read_master_translator:av_read
	wire   [63:0] msgdma_0_dma_read_master_readdata;                                                                  // mSGDMA_0_dma_read_master_translator:av_readdata -> mSGDMA_0:dma_read_master_readdata
	wire          msgdma_0_dma_read_master_readdatavalid;                                                             // mSGDMA_0_dma_read_master_translator:av_readdatavalid -> mSGDMA_0:dma_read_master_readdatavalid
	wire    [7:0] msgdma_0_dma_read_master_byteenable;                                                                // mSGDMA_0:dma_read_master_byteenable -> mSGDMA_0_dma_read_master_translator:av_byteenable
	wire    [5:0] msgdma_0_dma_write_master_burstcount;                                                               // mSGDMA_0:dma_write_master_burstcount -> mSGDMA_0_dma_write_master_translator:av_burstcount
	wire          msgdma_0_dma_write_master_waitrequest;                                                              // mSGDMA_0_dma_write_master_translator:av_waitrequest -> mSGDMA_0:dma_write_master_waitrequest
	wire   [63:0] msgdma_0_dma_write_master_writedata;                                                                // mSGDMA_0:dma_write_master_writedata -> mSGDMA_0_dma_write_master_translator:av_writedata
	wire   [31:0] msgdma_0_dma_write_master_address;                                                                  // mSGDMA_0:dma_write_master_address -> mSGDMA_0_dma_write_master_translator:av_address
	wire          msgdma_0_dma_write_master_write;                                                                    // mSGDMA_0:dma_write_master_write -> mSGDMA_0_dma_write_master_translator:av_write
	wire    [7:0] msgdma_0_dma_write_master_byteenable;                                                               // mSGDMA_0:dma_write_master_byteenable -> mSGDMA_0_dma_write_master_translator:av_byteenable
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_waitrequest;                                // mem_if_lpddr2_emif_0:avl_ready -> mem_if_lpddr2_emif_0_avl_translator:av_waitrequest
	wire   [10:0] mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_burstcount;                                 // mem_if_lpddr2_emif_0_avl_translator:av_burstcount -> mem_if_lpddr2_emif_0:avl_size
	wire   [63:0] mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_writedata;                                  // mem_if_lpddr2_emif_0_avl_translator:av_writedata -> mem_if_lpddr2_emif_0:avl_wdata
	wire   [23:0] mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_address;                                    // mem_if_lpddr2_emif_0_avl_translator:av_address -> mem_if_lpddr2_emif_0:avl_addr
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_write;                                      // mem_if_lpddr2_emif_0_avl_translator:av_write -> mem_if_lpddr2_emif_0:avl_write_req
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer;                         // mem_if_lpddr2_emif_0_avl_translator:av_beginbursttransfer -> mem_if_lpddr2_emif_0:avl_burstbegin
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_read;                                       // mem_if_lpddr2_emif_0_avl_translator:av_read -> mem_if_lpddr2_emif_0:avl_read_req
	wire   [63:0] mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdata;                                   // mem_if_lpddr2_emif_0:avl_rdata -> mem_if_lpddr2_emif_0_avl_translator:av_readdata
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid;                              // mem_if_lpddr2_emif_0:avl_rdata_valid -> mem_if_lpddr2_emif_0_avl_translator:av_readdatavalid
	wire    [7:0] mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_byteenable;                                 // mem_if_lpddr2_emif_0_avl_translator:av_byteenable -> mem_if_lpddr2_emif_0:avl_be
	wire          master_0_master_translator_avalon_universal_master_0_waitrequest;                                   // master_0_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_0_master_translator:uav_waitrequest
	wire    [2:0] master_0_master_translator_avalon_universal_master_0_burstcount;                                    // master_0_master_translator:uav_burstcount -> master_0_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_writedata;                                     // master_0_master_translator:uav_writedata -> master_0_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_address;                                       // master_0_master_translator:uav_address -> master_0_master_translator_avalon_universal_master_0_agent:av_address
	wire          master_0_master_translator_avalon_universal_master_0_lock;                                          // master_0_master_translator:uav_lock -> master_0_master_translator_avalon_universal_master_0_agent:av_lock
	wire          master_0_master_translator_avalon_universal_master_0_write;                                         // master_0_master_translator:uav_write -> master_0_master_translator_avalon_universal_master_0_agent:av_write
	wire          master_0_master_translator_avalon_universal_master_0_read;                                          // master_0_master_translator:uav_read -> master_0_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_readdata;                                      // master_0_master_translator_avalon_universal_master_0_agent:av_readdata -> master_0_master_translator:uav_readdata
	wire          master_0_master_translator_avalon_universal_master_0_debugaccess;                                   // master_0_master_translator:uav_debugaccess -> master_0_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] master_0_master_translator_avalon_universal_master_0_byteenable;                                    // master_0_master_translator:uav_byteenable -> master_0_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          master_0_master_translator_avalon_universal_master_0_readdatavalid;                                 // master_0_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_0_master_translator:uav_readdatavalid
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_waitrequest;              // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_driver_msgdma_0_avalon_master_translator:uav_waitrequest
	wire    [2:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_burstcount;               // master_driver_msgdma_0_avalon_master_translator:uav_burstcount -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_writedata;                // master_driver_msgdma_0_avalon_master_translator:uav_writedata -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_address;                  // master_driver_msgdma_0_avalon_master_translator:uav_address -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_lock;                     // master_driver_msgdma_0_avalon_master_translator:uav_lock -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_write;                    // master_driver_msgdma_0_avalon_master_translator:uav_write -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_read;                     // master_driver_msgdma_0_avalon_master_translator:uav_read -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdata;                 // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> master_driver_msgdma_0_avalon_master_translator:uav_readdata
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_debugaccess;              // master_driver_msgdma_0_avalon_master_translator:uav_debugaccess -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_byteenable;               // master_driver_msgdma_0_avalon_master_translator:uav_byteenable -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;            // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_driver_msgdma_0_avalon_master_translator:uav_readdatavalid
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // master_driver_msgdma_0_csr_translator:uav_waitrequest -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> master_driver_msgdma_0_csr_translator:uav_burstcount
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                  // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> master_driver_msgdma_0_csr_translator:uav_writedata
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_address;                    // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_address -> master_driver_msgdma_0_csr_translator:uav_address
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_write;                      // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_write -> master_driver_msgdma_0_csr_translator:uav_write
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_lock;                       // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_lock -> master_driver_msgdma_0_csr_translator:uav_lock
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_read;                       // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_read -> master_driver_msgdma_0_csr_translator:uav_read
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                   // master_driver_msgdma_0_csr_translator:uav_readdata -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // master_driver_msgdma_0_csr_translator:uav_readdatavalid -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> master_driver_msgdma_0_csr_translator:uav_debugaccess
	wire    [3:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> master_driver_msgdma_0_csr_translator:uav_byteenable
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;               // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;               // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // product_info_0_avalon_slave_0_translator:uav_waitrequest -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> product_info_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> product_info_0_avalon_slave_0_translator:uav_writedata
	wire   [31:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> product_info_0_avalon_slave_0_translator:uav_address
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> product_info_0_avalon_slave_0_translator:uav_write
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> product_info_0_avalon_slave_0_translator:uav_lock
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> product_info_0_avalon_slave_0_translator:uav_read
	wire   [31:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // product_info_0_avalon_slave_0_translator:uav_readdata -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // product_info_0_avalon_slave_0_translator:uav_readdatavalid -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> product_info_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> product_info_0_avalon_slave_0_translator:uav_byteenable
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // mSGDMA_0_mm_bridge_slv_translator:uav_waitrequest -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_burstcount -> mSGDMA_0_mm_bridge_slv_translator:uav_burstcount
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_writedata;                      // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_writedata -> mSGDMA_0_mm_bridge_slv_translator:uav_writedata
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_address;                        // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_address -> mSGDMA_0_mm_bridge_slv_translator:uav_address
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_write;                          // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_write -> mSGDMA_0_mm_bridge_slv_translator:uav_write
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_lock;                           // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_lock -> mSGDMA_0_mm_bridge_slv_translator:uav_lock
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_read;                           // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_read -> mSGDMA_0_mm_bridge_slv_translator:uav_read
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdata;                       // mSGDMA_0_mm_bridge_slv_translator:uav_readdata -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // mSGDMA_0_mm_bridge_slv_translator:uav_readdatavalid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mSGDMA_0_mm_bridge_slv_translator:uav_debugaccess
	wire    [3:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:m0_byteenable -> mSGDMA_0_mm_bridge_slv_translator:uav_byteenable
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_source_valid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_data;                    // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_source_data -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_waitrequest;                          // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> mSGDMA_0_dma_read_master_translator:uav_waitrequest
	wire    [8:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_burstcount;                           // mSGDMA_0_dma_read_master_translator:uav_burstcount -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_writedata;                            // mSGDMA_0_dma_read_master_translator:uav_writedata -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_address;                              // mSGDMA_0_dma_read_master_translator:uav_address -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_lock;                                 // mSGDMA_0_dma_read_master_translator:uav_lock -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_write;                                // mSGDMA_0_dma_read_master_translator:uav_write -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_read;                                 // mSGDMA_0_dma_read_master_translator:uav_read -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdata;                             // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> mSGDMA_0_dma_read_master_translator:uav_readdata
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_debugaccess;                          // mSGDMA_0_dma_read_master_translator:uav_debugaccess -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_byteenable;                           // mSGDMA_0_dma_read_master_translator:uav_byteenable -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdatavalid;                        // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> mSGDMA_0_dma_read_master_translator:uav_readdatavalid
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_waitrequest;                         // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> mSGDMA_0_dma_write_master_translator:uav_waitrequest
	wire    [8:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_burstcount;                          // mSGDMA_0_dma_write_master_translator:uav_burstcount -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_writedata;                           // mSGDMA_0_dma_write_master_translator:uav_writedata -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_address;                             // mSGDMA_0_dma_write_master_translator:uav_address -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_lock;                                // mSGDMA_0_dma_write_master_translator:uav_lock -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_write;                               // mSGDMA_0_dma_write_master_translator:uav_write -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_read;                                // mSGDMA_0_dma_write_master_translator:uav_read -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdata;                            // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> mSGDMA_0_dma_write_master_translator:uav_readdata
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_debugaccess;                         // mSGDMA_0_dma_write_master_translator:uav_debugaccess -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_byteenable;                          // mSGDMA_0_dma_write_master_translator:uav_byteenable -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdatavalid;                       // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> mSGDMA_0_dma_write_master_translator:uav_readdatavalid
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // mem_if_lpddr2_emif_0_avl_translator:uav_waitrequest -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [13:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> mem_if_lpddr2_emif_0_avl_translator:uav_burstcount
	wire   [63:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata;                    // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> mem_if_lpddr2_emif_0_avl_translator:uav_writedata
	wire   [31:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address;                      // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_address -> mem_if_lpddr2_emif_0_avl_translator:uav_address
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write;                        // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_write -> mem_if_lpddr2_emif_0_avl_translator:uav_write
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock;                         // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_lock -> mem_if_lpddr2_emif_0_avl_translator:uav_lock
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read;                         // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_read -> mem_if_lpddr2_emif_0_avl_translator:uav_read
	wire   [63:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                     // mem_if_lpddr2_emif_0_avl_translator:uav_readdata -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // mem_if_lpddr2_emif_0_avl_translator:uav_readdatavalid -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mem_if_lpddr2_emif_0_avl_translator:uav_debugaccess
	wire    [7:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> mem_if_lpddr2_emif_0_avl_translator:uav_byteenable
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [159:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data;                  // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [159:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [63:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // master_0_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_valid;                                // master_0_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // master_0_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [102:0] master_0_master_translator_avalon_universal_master_0_agent_cp_data;                                 // master_0_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router:sink_ready -> master_0_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;     // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;           // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;   // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [102:0] master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;            // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;           // addr_router_001:sink_ready -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                       // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [158:0] msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                        // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_002:sink_ready -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                      // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;              // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [158:0] msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                       // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_003:sink_ready -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [102:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire    [2:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> master_0_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> master_0_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> master_0_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                              // master_0_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mSGDMA_0:reset_reset_n]
	wire          master_driver_msgdma_0_reset_source_reset;                                                          // master_driver_msgdma_0:reset_out -> [rst_controller:reset_in0, rst_controller_005:reset_in0]
	wire          mem_if_lpddr2_emif_0_afi_reset_reset;                                                               // mem_if_lpddr2_emif_0:afi_reset_n -> [rst_controller:reset_in2, rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_005:reset_in2, rst_controller_006:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> mSGDMA_0:reset_0_reset_n
	wire          rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> [addr_router:reset, agent_pipeline_002:reset, agent_pipeline_003:reset, cmd_xbar_demux:reset, crosser:in_reset, crosser_002:out_reset, id_router_001:reset, limiter:reset, limiter_pipeline:reset, limiter_pipeline_001:reset, master_0_master_translator:reset, master_0_master_translator_avalon_universal_master_0_agent:reset, mux_pipeline_001:reset, mux_pipeline_004:reset, mux_pipeline_005:reset, mux_pipeline_006:reset, product_info_0:reset_n, product_info_0_avalon_slave_0_translator:reset, product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux:reset]
	wire          rst_controller_003_reset_out_reset;                                                                 // rst_controller_003:reset_out -> [addr_router_001:reset, agent_pipeline:reset, agent_pipeline_001:reset, cmd_xbar_demux_001:reset, crosser_001:in_reset, crosser_003:out_reset, id_router:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, master_driver_msgdma_0:reset_n, master_driver_msgdma_0_avalon_master_translator:reset, master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:reset, master_driver_msgdma_0_csr_translator:reset, master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:reset, master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mux_pipeline:reset, mux_pipeline_007:reset, rsp_xbar_demux:reset]
	wire          rst_controller_004_reset_out_reset;                                                                 // rst_controller_004:reset_out -> pll_0:rst
	wire          rst_controller_005_reset_out_reset;                                                                 // rst_controller_005:reset_out -> [addr_router_002:reset, addr_router_003:reset, agent_pipeline_004:reset, agent_pipeline_005:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux_002:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, id_router_002:reset, mSGDMA_0_dma_read_master_translator:reset, mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:reset, mSGDMA_0_dma_write_master_translator:reset, mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:reset, mSGDMA_0_mm_bridge_slv_translator:reset, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:reset, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mux_pipeline_002:reset, mux_pipeline_003:reset, mux_pipeline_010:reset, mux_pipeline_011:reset, rsp_xbar_demux_002:reset]
	wire          rst_controller_006_reset_out_reset;                                                                 // rst_controller_006:reset_out -> [agent_pipeline_006:reset, agent_pipeline_007:reset, cmd_xbar_mux_003:reset, id_router_003:reset, mem_if_lpddr2_emif_0_avl_translator:reset, mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:reset, mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mux_pipeline_008:reset, mux_pipeline_009:reset, rsp_xbar_demux_003:reset]
	wire          addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [102:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [2:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          mux_pipeline_007_source0_ready;                                                                     // master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> mux_pipeline_007:out_ready
	wire          id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [102:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [2:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [102:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [2:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [102:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [2:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [158:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [1:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          mux_pipeline_010_source0_ready;                                                                     // mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> mux_pipeline_010:out_ready
	wire          addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [158:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [1:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          mux_pipeline_011_source0_ready;                                                                     // mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> mux_pipeline_011:out_ready
	wire          id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [158:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [1:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> crosser:in_startofpacket
	wire  [102:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> crosser:in_data
	wire    [2:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                          // crosser:in_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> crosser_001:in_data
	wire    [2:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                      // crosser_001:in_ready -> cmd_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> crosser_002:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> crosser_002:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> crosser_002:in_data
	wire    [2:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> crosser_002:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                      // crosser_002:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                // rsp_xbar_demux_002:src1_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                      // rsp_xbar_demux_002:src1_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                              // rsp_xbar_demux_002:src1_startofpacket -> crosser_003:in_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src1_data;                                                                       // rsp_xbar_demux_002:src1_data -> crosser_003:in_data
	wire    [2:0] rsp_xbar_demux_002_src1_channel;                                                                    // rsp_xbar_demux_002:src1_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                      // crosser_003:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          limiter_pipeline_source0_endofpacket;                                                               // limiter_pipeline:out_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_pipeline_source0_valid;                                                                     // limiter_pipeline:out_valid -> cmd_xbar_demux:sink_valid
	wire          limiter_pipeline_source0_startofpacket;                                                             // limiter_pipeline:out_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [102:0] limiter_pipeline_source0_data;                                                                      // limiter_pipeline:out_data -> cmd_xbar_demux:sink_data
	wire    [2:0] limiter_pipeline_source0_channel;                                                                   // limiter_pipeline:out_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_pipeline_source0_ready;                                                                     // cmd_xbar_demux:sink_ready -> limiter_pipeline:out_ready
	wire          limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> limiter_pipeline:in_endofpacket
	wire    [0:0] limiter_cmd_src_valid;                                                                              // limiter:cmd_src_valid -> limiter_pipeline:in_valid
	wire          limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> limiter_pipeline:in_startofpacket
	wire  [102:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> limiter_pipeline:in_data
	wire    [2:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> limiter_pipeline:in_channel
	wire          limiter_cmd_src_ready;                                                                              // limiter_pipeline:in_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter_pipeline_001:in_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter_pipeline_001:in_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter_pipeline_001:in_startofpacket
	wire  [102:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter_pipeline_001:in_data
	wire    [2:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter_pipeline_001:in_channel
	wire          rsp_xbar_mux_src_ready;                                                                             // limiter_pipeline_001:in_ready -> rsp_xbar_mux:src_ready
	wire          limiter_pipeline_001_source0_endofpacket;                                                           // limiter_pipeline_001:out_endofpacket -> limiter:rsp_sink_endofpacket
	wire          limiter_pipeline_001_source0_valid;                                                                 // limiter_pipeline_001:out_valid -> limiter:rsp_sink_valid
	wire          limiter_pipeline_001_source0_startofpacket;                                                         // limiter_pipeline_001:out_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [102:0] limiter_pipeline_001_source0_data;                                                                  // limiter_pipeline_001:out_data -> limiter:rsp_sink_data
	wire    [2:0] limiter_pipeline_001_source0_channel;                                                               // limiter_pipeline_001:out_channel -> limiter:rsp_sink_channel
	wire          limiter_pipeline_001_source0_ready;                                                                 // limiter:rsp_sink_ready -> limiter_pipeline_001:out_ready
	wire          mux_pipeline_source0_ready;                                                                         // agent_pipeline:in_ready -> mux_pipeline:out_ready
	wire          agent_pipeline_source0_endofpacket;                                                                 // agent_pipeline:out_endofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_source0_valid;                                                                       // agent_pipeline:out_valid -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_source0_startofpacket;                                                               // agent_pipeline:out_startofpacket -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] agent_pipeline_source0_data;                                                                        // agent_pipeline:out_data -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] agent_pipeline_source0_channel;                                                                     // agent_pipeline:out_channel -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_source0_ready;                                                                       // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline:out_ready
	wire          agent_pipeline_001_source0_endofpacket;                                                             // agent_pipeline_001:out_endofpacket -> id_router:sink_endofpacket
	wire          agent_pipeline_001_source0_valid;                                                                   // agent_pipeline_001:out_valid -> id_router:sink_valid
	wire          agent_pipeline_001_source0_startofpacket;                                                           // agent_pipeline_001:out_startofpacket -> id_router:sink_startofpacket
	wire  [102:0] agent_pipeline_001_source0_data;                                                                    // agent_pipeline_001:out_data -> id_router:sink_data
	wire          agent_pipeline_001_source0_ready;                                                                   // id_router:sink_ready -> agent_pipeline_001:out_ready
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_001:in_endofpacket
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_valid;                      // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_001:in_valid
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_001:in_startofpacket
	wire  [102:0] master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_data;                       // master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_001:in_data
	wire          master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_ready;                      // agent_pipeline_001:in_ready -> master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_001_source0_ready;                                                                     // agent_pipeline_002:in_ready -> mux_pipeline_001:out_ready
	wire          agent_pipeline_002_source0_endofpacket;                                                             // agent_pipeline_002:out_endofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_002_source0_valid;                                                                   // agent_pipeline_002:out_valid -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_002_source0_startofpacket;                                                           // agent_pipeline_002:out_startofpacket -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] agent_pipeline_002_source0_data;                                                                    // agent_pipeline_002:out_data -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] agent_pipeline_002_source0_channel;                                                                 // agent_pipeline_002:out_channel -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_002_source0_ready;                                                                   // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_002:out_ready
	wire          agent_pipeline_003_source0_endofpacket;                                                             // agent_pipeline_003:out_endofpacket -> id_router_001:sink_endofpacket
	wire          agent_pipeline_003_source0_valid;                                                                   // agent_pipeline_003:out_valid -> id_router_001:sink_valid
	wire          agent_pipeline_003_source0_startofpacket;                                                           // agent_pipeline_003:out_startofpacket -> id_router_001:sink_startofpacket
	wire  [102:0] agent_pipeline_003_source0_data;                                                                    // agent_pipeline_003:out_data -> id_router_001:sink_data
	wire          agent_pipeline_003_source0_ready;                                                                   // id_router_001:sink_ready -> agent_pipeline_003:out_ready
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_003:in_endofpacket
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_003:in_valid
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_003:in_startofpacket
	wire  [102:0] product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_003:in_data
	wire          product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // agent_pipeline_003:in_ready -> product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                   // cmd_xbar_mux_002:src_endofpacket -> agent_pipeline_004:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                         // cmd_xbar_mux_002:src_valid -> agent_pipeline_004:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                 // cmd_xbar_mux_002:src_startofpacket -> agent_pipeline_004:in_startofpacket
	wire  [102:0] cmd_xbar_mux_002_src_data;                                                                          // cmd_xbar_mux_002:src_data -> agent_pipeline_004:in_data
	wire    [2:0] cmd_xbar_mux_002_src_channel;                                                                       // cmd_xbar_mux_002:src_channel -> agent_pipeline_004:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                         // agent_pipeline_004:in_ready -> cmd_xbar_mux_002:src_ready
	wire          agent_pipeline_004_source0_endofpacket;                                                             // agent_pipeline_004:out_endofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_004_source0_valid;                                                                   // agent_pipeline_004:out_valid -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_004_source0_startofpacket;                                                           // agent_pipeline_004:out_startofpacket -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] agent_pipeline_004_source0_data;                                                                    // agent_pipeline_004:out_data -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] agent_pipeline_004_source0_channel;                                                                 // agent_pipeline_004:out_channel -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_004_source0_ready;                                                                   // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_004:out_ready
	wire          agent_pipeline_005_source0_endofpacket;                                                             // agent_pipeline_005:out_endofpacket -> id_router_002:sink_endofpacket
	wire          agent_pipeline_005_source0_valid;                                                                   // agent_pipeline_005:out_valid -> id_router_002:sink_valid
	wire          agent_pipeline_005_source0_startofpacket;                                                           // agent_pipeline_005:out_startofpacket -> id_router_002:sink_startofpacket
	wire  [102:0] agent_pipeline_005_source0_data;                                                                    // agent_pipeline_005:out_data -> id_router_002:sink_data
	wire          agent_pipeline_005_source0_ready;                                                                   // id_router_002:sink_ready -> agent_pipeline_005:out_ready
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_005:in_endofpacket
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_valid;                          // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_005:in_valid
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_005:in_startofpacket
	wire  [102:0] msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_data;                           // mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_005:in_data
	wire          msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_ready;                          // agent_pipeline_005:in_ready -> mSGDMA_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                   // cmd_xbar_mux_003:src_endofpacket -> agent_pipeline_006:in_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                         // cmd_xbar_mux_003:src_valid -> agent_pipeline_006:in_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                 // cmd_xbar_mux_003:src_startofpacket -> agent_pipeline_006:in_startofpacket
	wire  [158:0] cmd_xbar_mux_003_src_data;                                                                          // cmd_xbar_mux_003:src_data -> agent_pipeline_006:in_data
	wire    [1:0] cmd_xbar_mux_003_src_channel;                                                                       // cmd_xbar_mux_003:src_channel -> agent_pipeline_006:in_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                         // agent_pipeline_006:in_ready -> cmd_xbar_mux_003:src_ready
	wire          agent_pipeline_006_source0_endofpacket;                                                             // agent_pipeline_006:out_endofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_006_source0_valid;                                                                   // agent_pipeline_006:out_valid -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_006_source0_startofpacket;                                                           // agent_pipeline_006:out_startofpacket -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [158:0] agent_pipeline_006_source0_data;                                                                    // agent_pipeline_006:out_data -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] agent_pipeline_006_source0_channel;                                                                 // agent_pipeline_006:out_channel -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_006_source0_ready;                                                                   // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_006:out_ready
	wire          agent_pipeline_007_source0_endofpacket;                                                             // agent_pipeline_007:out_endofpacket -> id_router_003:sink_endofpacket
	wire          agent_pipeline_007_source0_valid;                                                                   // agent_pipeline_007:out_valid -> id_router_003:sink_valid
	wire          agent_pipeline_007_source0_startofpacket;                                                           // agent_pipeline_007:out_startofpacket -> id_router_003:sink_startofpacket
	wire  [158:0] agent_pipeline_007_source0_data;                                                                    // agent_pipeline_007:out_data -> id_router_003:sink_data
	wire          agent_pipeline_007_source0_ready;                                                                   // id_router_003:sink_ready -> agent_pipeline_007:out_ready
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_007:in_endofpacket
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid;                        // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_007:in_valid
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_007:in_startofpacket
	wire  [158:0] mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data;                         // mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_007:in_data
	wire          mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready;                        // agent_pipeline_007:in_ready -> mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> mux_pipeline:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> mux_pipeline:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> mux_pipeline:in_startofpacket
	wire  [102:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> mux_pipeline:in_data
	wire    [2:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> mux_pipeline:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                                          // mux_pipeline:in_ready -> cmd_xbar_demux:src0_ready
	wire          mux_pipeline_source0_endofpacket;                                                                   // mux_pipeline:out_endofpacket -> agent_pipeline:in_endofpacket
	wire          mux_pipeline_source0_valid;                                                                         // mux_pipeline:out_valid -> agent_pipeline:in_valid
	wire          mux_pipeline_source0_startofpacket;                                                                 // mux_pipeline:out_startofpacket -> agent_pipeline:in_startofpacket
	wire  [102:0] mux_pipeline_source0_data;                                                                          // mux_pipeline:out_data -> agent_pipeline:in_data
	wire    [2:0] mux_pipeline_source0_channel;                                                                       // mux_pipeline:out_channel -> agent_pipeline:in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> mux_pipeline_001:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> mux_pipeline_001:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> mux_pipeline_001:in_startofpacket
	wire  [102:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> mux_pipeline_001:in_data
	wire    [2:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> mux_pipeline_001:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                          // mux_pipeline_001:in_ready -> cmd_xbar_demux:src1_ready
	wire          mux_pipeline_001_source0_endofpacket;                                                               // mux_pipeline_001:out_endofpacket -> agent_pipeline_002:in_endofpacket
	wire          mux_pipeline_001_source0_valid;                                                                     // mux_pipeline_001:out_valid -> agent_pipeline_002:in_valid
	wire          mux_pipeline_001_source0_startofpacket;                                                             // mux_pipeline_001:out_startofpacket -> agent_pipeline_002:in_startofpacket
	wire  [102:0] mux_pipeline_001_source0_data;                                                                      // mux_pipeline_001:out_data -> agent_pipeline_002:in_data
	wire    [2:0] mux_pipeline_001_source0_channel;                                                                   // mux_pipeline_001:out_channel -> agent_pipeline_002:in_channel
	wire          crosser_out_endofpacket;                                                                            // crosser:out_endofpacket -> mux_pipeline_002:in_endofpacket
	wire          crosser_out_valid;                                                                                  // crosser:out_valid -> mux_pipeline_002:in_valid
	wire          crosser_out_startofpacket;                                                                          // crosser:out_startofpacket -> mux_pipeline_002:in_startofpacket
	wire  [102:0] crosser_out_data;                                                                                   // crosser:out_data -> mux_pipeline_002:in_data
	wire    [2:0] crosser_out_channel;                                                                                // crosser:out_channel -> mux_pipeline_002:in_channel
	wire          crosser_out_ready;                                                                                  // mux_pipeline_002:in_ready -> crosser:out_ready
	wire          mux_pipeline_002_source0_endofpacket;                                                               // mux_pipeline_002:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          mux_pipeline_002_source0_valid;                                                                     // mux_pipeline_002:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          mux_pipeline_002_source0_startofpacket;                                                             // mux_pipeline_002:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [102:0] mux_pipeline_002_source0_data;                                                                      // mux_pipeline_002:out_data -> cmd_xbar_mux_002:sink0_data
	wire    [2:0] mux_pipeline_002_source0_channel;                                                                   // mux_pipeline_002:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          mux_pipeline_002_source0_ready;                                                                     // cmd_xbar_mux_002:sink0_ready -> mux_pipeline_002:out_ready
	wire          crosser_001_out_endofpacket;                                                                        // crosser_001:out_endofpacket -> mux_pipeline_003:in_endofpacket
	wire          crosser_001_out_valid;                                                                              // crosser_001:out_valid -> mux_pipeline_003:in_valid
	wire          crosser_001_out_startofpacket;                                                                      // crosser_001:out_startofpacket -> mux_pipeline_003:in_startofpacket
	wire  [102:0] crosser_001_out_data;                                                                               // crosser_001:out_data -> mux_pipeline_003:in_data
	wire    [2:0] crosser_001_out_channel;                                                                            // crosser_001:out_channel -> mux_pipeline_003:in_channel
	wire          crosser_001_out_ready;                                                                              // mux_pipeline_003:in_ready -> crosser_001:out_ready
	wire          mux_pipeline_003_source0_endofpacket;                                                               // mux_pipeline_003:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          mux_pipeline_003_source0_valid;                                                                     // mux_pipeline_003:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          mux_pipeline_003_source0_startofpacket;                                                             // mux_pipeline_003:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [102:0] mux_pipeline_003_source0_data;                                                                      // mux_pipeline_003:out_data -> cmd_xbar_mux_002:sink1_data
	wire    [2:0] mux_pipeline_003_source0_channel;                                                                   // mux_pipeline_003:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          mux_pipeline_003_source0_ready;                                                                     // cmd_xbar_mux_002:sink1_ready -> mux_pipeline_003:out_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> mux_pipeline_004:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> mux_pipeline_004:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> mux_pipeline_004:in_startofpacket
	wire  [102:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> mux_pipeline_004:in_data
	wire    [2:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> mux_pipeline_004:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                                          // mux_pipeline_004:in_ready -> rsp_xbar_demux:src0_ready
	wire          mux_pipeline_004_source0_endofpacket;                                                               // mux_pipeline_004:out_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          mux_pipeline_004_source0_valid;                                                                     // mux_pipeline_004:out_valid -> rsp_xbar_mux:sink0_valid
	wire          mux_pipeline_004_source0_startofpacket;                                                             // mux_pipeline_004:out_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [102:0] mux_pipeline_004_source0_data;                                                                      // mux_pipeline_004:out_data -> rsp_xbar_mux:sink0_data
	wire    [2:0] mux_pipeline_004_source0_channel;                                                                   // mux_pipeline_004:out_channel -> rsp_xbar_mux:sink0_channel
	wire          mux_pipeline_004_source0_ready;                                                                     // rsp_xbar_mux:sink0_ready -> mux_pipeline_004:out_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> mux_pipeline_005:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> mux_pipeline_005:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> mux_pipeline_005:in_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> mux_pipeline_005:in_data
	wire    [2:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> mux_pipeline_005:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                      // mux_pipeline_005:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          mux_pipeline_005_source0_endofpacket;                                                               // mux_pipeline_005:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          mux_pipeline_005_source0_valid;                                                                     // mux_pipeline_005:out_valid -> rsp_xbar_mux:sink1_valid
	wire          mux_pipeline_005_source0_startofpacket;                                                             // mux_pipeline_005:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [102:0] mux_pipeline_005_source0_data;                                                                      // mux_pipeline_005:out_data -> rsp_xbar_mux:sink1_data
	wire    [2:0] mux_pipeline_005_source0_channel;                                                                   // mux_pipeline_005:out_channel -> rsp_xbar_mux:sink1_channel
	wire          mux_pipeline_005_source0_ready;                                                                     // rsp_xbar_mux:sink1_ready -> mux_pipeline_005:out_ready
	wire          crosser_002_out_endofpacket;                                                                        // crosser_002:out_endofpacket -> mux_pipeline_006:in_endofpacket
	wire          crosser_002_out_valid;                                                                              // crosser_002:out_valid -> mux_pipeline_006:in_valid
	wire          crosser_002_out_startofpacket;                                                                      // crosser_002:out_startofpacket -> mux_pipeline_006:in_startofpacket
	wire  [102:0] crosser_002_out_data;                                                                               // crosser_002:out_data -> mux_pipeline_006:in_data
	wire    [2:0] crosser_002_out_channel;                                                                            // crosser_002:out_channel -> mux_pipeline_006:in_channel
	wire          crosser_002_out_ready;                                                                              // mux_pipeline_006:in_ready -> crosser_002:out_ready
	wire          mux_pipeline_006_source0_endofpacket;                                                               // mux_pipeline_006:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          mux_pipeline_006_source0_valid;                                                                     // mux_pipeline_006:out_valid -> rsp_xbar_mux:sink2_valid
	wire          mux_pipeline_006_source0_startofpacket;                                                             // mux_pipeline_006:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [102:0] mux_pipeline_006_source0_data;                                                                      // mux_pipeline_006:out_data -> rsp_xbar_mux:sink2_data
	wire    [2:0] mux_pipeline_006_source0_channel;                                                                   // mux_pipeline_006:out_channel -> rsp_xbar_mux:sink2_channel
	wire          mux_pipeline_006_source0_ready;                                                                     // rsp_xbar_mux:sink2_ready -> mux_pipeline_006:out_ready
	wire          crosser_003_out_endofpacket;                                                                        // crosser_003:out_endofpacket -> mux_pipeline_007:in_endofpacket
	wire          crosser_003_out_valid;                                                                              // crosser_003:out_valid -> mux_pipeline_007:in_valid
	wire          crosser_003_out_startofpacket;                                                                      // crosser_003:out_startofpacket -> mux_pipeline_007:in_startofpacket
	wire  [102:0] crosser_003_out_data;                                                                               // crosser_003:out_data -> mux_pipeline_007:in_data
	wire    [2:0] crosser_003_out_channel;                                                                            // crosser_003:out_channel -> mux_pipeline_007:in_channel
	wire          crosser_003_out_ready;                                                                              // mux_pipeline_007:in_ready -> crosser_003:out_ready
	wire          mux_pipeline_007_source0_endofpacket;                                                               // mux_pipeline_007:out_endofpacket -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          mux_pipeline_007_source0_valid;                                                                     // mux_pipeline_007:out_valid -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          mux_pipeline_007_source0_startofpacket;                                                             // mux_pipeline_007:out_startofpacket -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] mux_pipeline_007_source0_data;                                                                      // mux_pipeline_007:out_data -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] mux_pipeline_007_source0_channel;                                                                   // mux_pipeline_007:out_channel -> master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> mux_pipeline_008:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> mux_pipeline_008:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> mux_pipeline_008:in_startofpacket
	wire  [158:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> mux_pipeline_008:in_data
	wire    [1:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> mux_pipeline_008:in_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                      // mux_pipeline_008:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          mux_pipeline_008_source0_endofpacket;                                                               // mux_pipeline_008:out_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          mux_pipeline_008_source0_valid;                                                                     // mux_pipeline_008:out_valid -> cmd_xbar_mux_003:sink0_valid
	wire          mux_pipeline_008_source0_startofpacket;                                                             // mux_pipeline_008:out_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [158:0] mux_pipeline_008_source0_data;                                                                      // mux_pipeline_008:out_data -> cmd_xbar_mux_003:sink0_data
	wire    [1:0] mux_pipeline_008_source0_channel;                                                                   // mux_pipeline_008:out_channel -> cmd_xbar_mux_003:sink0_channel
	wire          mux_pipeline_008_source0_ready;                                                                     // cmd_xbar_mux_003:sink0_ready -> mux_pipeline_008:out_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> mux_pipeline_009:in_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> mux_pipeline_009:in_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> mux_pipeline_009:in_startofpacket
	wire  [158:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> mux_pipeline_009:in_data
	wire    [1:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> mux_pipeline_009:in_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                      // mux_pipeline_009:in_ready -> cmd_xbar_demux_003:src0_ready
	wire          mux_pipeline_009_source0_endofpacket;                                                               // mux_pipeline_009:out_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          mux_pipeline_009_source0_valid;                                                                     // mux_pipeline_009:out_valid -> cmd_xbar_mux_003:sink1_valid
	wire          mux_pipeline_009_source0_startofpacket;                                                             // mux_pipeline_009:out_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [158:0] mux_pipeline_009_source0_data;                                                                      // mux_pipeline_009:out_data -> cmd_xbar_mux_003:sink1_data
	wire    [1:0] mux_pipeline_009_source0_channel;                                                                   // mux_pipeline_009:out_channel -> cmd_xbar_mux_003:sink1_channel
	wire          mux_pipeline_009_source0_ready;                                                                     // cmd_xbar_mux_003:sink1_ready -> mux_pipeline_009:out_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> mux_pipeline_010:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> mux_pipeline_010:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> mux_pipeline_010:in_startofpacket
	wire  [158:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> mux_pipeline_010:in_data
	wire    [1:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> mux_pipeline_010:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                      // mux_pipeline_010:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          mux_pipeline_010_source0_endofpacket;                                                               // mux_pipeline_010:out_endofpacket -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          mux_pipeline_010_source0_valid;                                                                     // mux_pipeline_010:out_valid -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          mux_pipeline_010_source0_startofpacket;                                                             // mux_pipeline_010:out_startofpacket -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [158:0] mux_pipeline_010_source0_data;                                                                      // mux_pipeline_010:out_data -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] mux_pipeline_010_source0_channel;                                                                   // mux_pipeline_010:out_channel -> mSGDMA_0_dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                // rsp_xbar_demux_003:src1_endofpacket -> mux_pipeline_011:in_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                      // rsp_xbar_demux_003:src1_valid -> mux_pipeline_011:in_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                              // rsp_xbar_demux_003:src1_startofpacket -> mux_pipeline_011:in_startofpacket
	wire  [158:0] rsp_xbar_demux_003_src1_data;                                                                       // rsp_xbar_demux_003:src1_data -> mux_pipeline_011:in_data
	wire    [1:0] rsp_xbar_demux_003_src1_channel;                                                                    // rsp_xbar_demux_003:src1_channel -> mux_pipeline_011:in_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                      // mux_pipeline_011:in_ready -> rsp_xbar_demux_003:src1_ready
	wire          mux_pipeline_011_source0_endofpacket;                                                               // mux_pipeline_011:out_endofpacket -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          mux_pipeline_011_source0_valid;                                                                     // mux_pipeline_011:out_valid -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          mux_pipeline_011_source0_startofpacket;                                                             // mux_pipeline_011:out_startofpacket -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [158:0] mux_pipeline_011_source0_data;                                                                      // mux_pipeline_011:out_data -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] mux_pipeline_011_source0_channel;                                                                   // mux_pipeline_011:out_channel -> mSGDMA_0_dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire    [1:0] master_driver_msgdma_0_interrupt_receiver_irq;                                                      // irq_mapper:sender_irq -> master_driver_msgdma_0:irq
	wire          irq_mapper_receiver0_irq;                                                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                      // mSGDMA_0:dispatcher_write_csr_irq_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                           // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                  // mSGDMA_0:dispatcher_read_csr_irq_irq -> irq_synchronizer_001:receiver_irq

	q_sys_mSGDMA_0 msgdma_0 (
		.mm_bridge_slv_waitrequest       (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_waitrequest),   //            mm_bridge_slv.waitrequest
		.mm_bridge_slv_readdata          (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdata),      //                         .readdata
		.mm_bridge_slv_readdatavalid     (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdatavalid), //                         .readdatavalid
		.mm_bridge_slv_burstcount        (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_burstcount),    //                         .burstcount
		.mm_bridge_slv_writedata         (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_writedata),     //                         .writedata
		.mm_bridge_slv_address           (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_address),       //                         .address
		.mm_bridge_slv_write             (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_write),         //                         .write
		.mm_bridge_slv_read              (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_read),          //                         .read
		.mm_bridge_slv_byteenable        (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_byteenable),    //                         .byteenable
		.mm_bridge_slv_debugaccess       (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_debugaccess),   //                         .debugaccess
		.reset_reset_n                   (~rst_controller_reset_out_reset),                                     //                    reset.reset_n
		.clk_clk                         (mem_if_lpddr2_emif_0_afi_clk_clk),                                    //                      clk.clk
		.dma_read_master_address         (msgdma_0_dma_read_master_address),                                    //          dma_read_master.address
		.dma_read_master_read            (msgdma_0_dma_read_master_read),                                       //                         .read
		.dma_read_master_byteenable      (msgdma_0_dma_read_master_byteenable),                                 //                         .byteenable
		.dma_read_master_readdata        (msgdma_0_dma_read_master_readdata),                                   //                         .readdata
		.dma_read_master_waitrequest     (msgdma_0_dma_read_master_waitrequest),                                //                         .waitrequest
		.dma_read_master_readdatavalid   (msgdma_0_dma_read_master_readdatavalid),                              //                         .readdatavalid
		.dma_read_master_burstcount      (msgdma_0_dma_read_master_burstcount),                                 //                         .burstcount
		.dma_write_master_address        (msgdma_0_dma_write_master_address),                                   //         dma_write_master.address
		.dma_write_master_write          (msgdma_0_dma_write_master_write),                                     //                         .write
		.dma_write_master_byteenable     (msgdma_0_dma_write_master_byteenable),                                //                         .byteenable
		.dma_write_master_writedata      (msgdma_0_dma_write_master_writedata),                                 //                         .writedata
		.dma_write_master_waitrequest    (msgdma_0_dma_write_master_waitrequest),                               //                         .waitrequest
		.dma_write_master_burstcount     (msgdma_0_dma_write_master_burstcount),                                //                         .burstcount
		.dispatcher_write_csr_irq_irq    (irq_synchronizer_receiver_irq),                                       // dispatcher_write_csr_irq.irq
		.dispatcher_read_csr_irq_irq     (irq_synchronizer_001_receiver_irq),                                   //  dispatcher_read_csr_irq.irq
		.clk_0_clk                       (clk_50_clk),                                                          //                    clk_0.clk
		.reset_0_reset_n                 (~rst_controller_001_reset_out_reset),                                 //                  reset_0.reset_n
		.status_mon_out_cal_fail_mon     (msgdma_0_status_mon_out_cal_fail_mon),                                //           status_mon_out.cal_fail_mon
		.status_mon_out_cal_success_mon  (msgdma_0_status_mon_out_cal_success_mon),                             //                         .cal_success_mon
		.status_mon_out_init_done_mon    (msgdma_0_status_mon_out_init_done_mon),                               //                         .init_done_mon
		.status_mon_in_local_init_done   (mem_if_lpddr2_emif_0_status_local_init_done),                         //            status_mon_in.local_init_done
		.status_mon_in_local_cal_success (mem_if_lpddr2_emif_0_status_local_cal_success),                       //                         .local_cal_success
		.status_mon_in_local_cal_fail    (mem_if_lpddr2_emif_0_status_local_cal_fail),                          //                         .local_cal_fail
		.reset_source_reset_n            ()                                                                     //             reset_source.reset_n
	);

	product_info product_info_0 (
		.clk          (clk_50_clk),                                                               //       clock_reset.clk
		.reset_n      (~rst_controller_002_reset_out_reset),                                      // clock_reset_reset.reset_n
		.chipselect_n (~product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //    avalon_slave_0.chipselect_n
		.read_n       (~product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_data_read (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_address   (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_address)      //                  .address
	);

	master_driver_msgdma #(
		.PRBS_PATTERN_GENERATOR_BASE (32'b00000000001000000000000001000000),
		.PRBS_PATTERN_CHECKER_BASE   (32'b00000000001000000000000000000000),
		.MEMORY_BASE_ADDRESS         (32'b00000000000000000000000000000000),
		.MEMORY_SPAN                 (32'b00001000000000000000000000000000),
		.BLOCK_SIZE                  (32'b00100000000000000000000000000000),
		.DISPATCHER_WRITE_CSR        (32'b00000000001000000000000001100000),
		.DISPATCHER_WRITE_DESCRIPTOR (32'b00000000001000000000000010100000),
		.DISPATCHER_READ_CSR         (32'b00000000001000000000000010000000),
		.DISPATCHER_READ_DESCRIPTOR  (32'b00000000001000000000000010110000),
		.TIMER_BASE                  (32'b00000000001010000001000000000000),
		.FREQUENCY_COUNTER_BASE      (32'b00000000001010010000000000000000),
		.ENABLE_PER_INFO             (1),
		.LOCAL_DATA_WORDS            (32'b00000000000000000000000000001000)
	) master_driver_msgdma_0 (
		.reset_n         (~rst_controller_003_reset_out_reset),                                   //              reset.reset_n
		.clk             (clk_50_clk),                                                            //              clock.clk
		.csr_address     (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_address),     //                csr.address
		.csr_read        (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_read),        //                   .read
		.csr_write       (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_write),       //                   .write
		.csr_readdata    (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.csr_writedata   (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.csr_waitrequest (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq             (master_driver_msgdma_0_interrupt_receiver_irq),                         // interrupt_receiver.irq
		.waitrequest_in  (master_driver_msgdma_0_avalon_master_waitrequest),                      //      avalon_master.waitrequest
		.csn             (master_driver_msgdma_0_avalon_master_chipselect),                       //                   .chipselect_n
		.wen             (master_driver_msgdma_0_avalon_master_write),                            //                   .write_n
		.oen             (master_driver_msgdma_0_avalon_master_read),                             //                   .read_n
		.be              (master_driver_msgdma_0_avalon_master_byteenable),                       //                   .byteenable
		.address         (master_driver_msgdma_0_avalon_master_address),                          //                   .address
		.data_write      (master_driver_msgdma_0_avalon_master_writedata),                        //                   .writedata
		.data_read       (master_driver_msgdma_0_avalon_master_readdata),                         //                   .readdata
		.reset_out       (master_driver_msgdma_0_reset_source_reset),                             //       reset_source.reset
		.error_mon       (master_driver_msgdma_0_conduit_end_error_mon),                          //        conduit_end.export
		.status_mon      (master_driver_msgdma_0_conduit_end_status_mon)                          //                   .export
	);

	q_sys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_50_clk),                    //          clk.clk
		.clk_reset_reset      (~reset_50_reset_n),             //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	q_sys_pll_0 pll_0 (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_004_reset_out_reset), //   reset.reset
		.outclk_0 (),                                   // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	q_sys_mem_if_lpddr2_emif_0 mem_if_lpddr2_emif_0 (
		.pll_ref_clk       (clk_clk),                                                                    //  pll_ref_clk.clk
		.global_reset_n    (reset_reset_n),                                                              // global_reset.reset_n
		.soft_reset_n      (reset_reset_n),                                                              //   soft_reset.reset_n
		.afi_clk           (mem_if_lpddr2_emif_0_afi_clk_clk),                                           //      afi_clk.clk
		.afi_half_clk      (),                                                                           // afi_half_clk.clk
		.afi_reset_n       (mem_if_lpddr2_emif_0_afi_reset_reset),                                       //    afi_reset.reset_n
		.mem_ca            (memory_mem_ca),                                                              //       memory.mem_ca
		.mem_ck            (memory_mem_ck),                                                              //             .mem_ck
		.mem_ck_n          (memory_mem_ck_n),                                                            //             .mem_ck_n
		.mem_cke           (memory_mem_cke),                                                             //             .mem_cke
		.mem_cs_n          (memory_mem_cs_n),                                                            //             .mem_cs_n
		.mem_dm            (memory_mem_dm),                                                              //             .mem_dm
		.mem_dq            (memory_mem_dq),                                                              //             .mem_dq
		.mem_dqs           (memory_mem_dqs),                                                             //             .mem_dqs
		.mem_dqs_n         (memory_mem_dqs_n),                                                           //             .mem_dqs_n
		.avl_ready         (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),        //          avl.waitrequest_n
		.avl_burstbegin    (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer), //             .beginbursttransfer
		.avl_addr          (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_address),            //             .address
		.avl_rdata_valid   (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),      //             .readdatavalid
		.avl_rdata         (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdata),           //             .readdata
		.avl_wdata         (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_writedata),          //             .writedata
		.avl_be            (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_byteenable),         //             .byteenable
		.avl_read_req      (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_read),               //             .read
		.avl_write_req     (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_write),              //             .write
		.avl_size          (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_burstcount),         //             .burstcount
		.local_init_done   (mem_if_lpddr2_emif_0_status_local_init_done),                                //       status.local_init_done
		.local_cal_success (mem_if_lpddr2_emif_0_status_local_cal_success),                              //             .local_cal_success
		.local_cal_fail    (mem_if_lpddr2_emif_0_status_local_cal_fail),                                 //             .local_cal_fail
		.oct_rzqin         (oct_rzqin)                                                                   //          oct.rzqin
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_0_master_translator (
		.clk                   (clk_50_clk),                                                         //                       clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                 //                     reset.reset
		.uav_address           (master_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (master_0_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (master_0_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (master_0_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (master_0_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (master_0_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (master_0_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (master_0_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (master_0_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (master_0_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (master_0_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (master_0_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (master_0_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (master_0_master_byteenable),                                         //                          .byteenable
		.av_read               (master_0_master_read),                                               //                          .read
		.av_readdata           (master_0_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (master_0_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (master_0_master_write),                                              //                          .write
		.av_writedata          (master_0_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_driver_msgdma_0_avalon_master_translator (
		.clk                   (clk_50_clk),                                                                              //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                      //                     reset.reset
		.uav_address           (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (master_driver_msgdma_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (master_driver_msgdma_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (master_driver_msgdma_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_chipselect         (~master_driver_msgdma_0_avalon_master_chipselect),                                        //                          .chipselect
		.av_read               (~master_driver_msgdma_0_avalon_master_read),                                              //                          .read
		.av_readdata           (master_driver_msgdma_0_avalon_master_readdata),                                           //                          .readdata
		.av_write              (~master_driver_msgdma_0_avalon_master_write),                                             //                          .write
		.av_writedata          (master_driver_msgdma_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                                    //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                                        //               (terminated)
		.av_lock               (1'b0),                                                                                    //               (terminated)
		.av_debugaccess        (1'b0),                                                                                    //               (terminated)
		.uav_clken             (),                                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                                     //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) master_driver_msgdma_0_csr_translator (
		.clk                   (clk_50_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (master_driver_msgdma_0_csr_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) product_info_0_avalon_slave_0_translator (
		.clk                   (clk_50_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_chipselect         (product_info_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_write              (),                                                                                         //              (terminated)
		.av_writedata          (),                                                                                         //              (terminated)
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) msgdma_0_mm_bridge_slv_translator (
		.clk                   (mem_if_lpddr2_emif_0_afi_clk_clk),                                                  //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                                //                    reset.reset
		.uav_address           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (msgdma_0_mm_bridge_slv_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (6),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (9),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) msgdma_0_dma_read_master_translator (
		.clk                   (mem_if_lpddr2_emif_0_afi_clk_clk),                                            //                       clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                          //                     reset.reset
		.uav_address           (msgdma_0_dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (msgdma_0_dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (msgdma_0_dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (msgdma_0_dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (msgdma_0_dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (msgdma_0_dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (msgdma_0_dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (msgdma_0_dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (msgdma_0_dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (msgdma_0_dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (msgdma_0_dma_read_master_burstcount),                                         //                          .burstcount
		.av_byteenable         (msgdma_0_dma_read_master_byteenable),                                         //                          .byteenable
		.av_read               (msgdma_0_dma_read_master_read),                                               //                          .read
		.av_readdata           (msgdma_0_dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (msgdma_0_dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (64'b0000000000000000000000000000000000000000000000000000000000000000),        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (6),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (9),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) msgdma_0_dma_write_master_translator (
		.clk                   (mem_if_lpddr2_emif_0_afi_clk_clk),                                             //                       clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                           //                     reset.reset
		.uav_address           (msgdma_0_dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (msgdma_0_dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (msgdma_0_dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (msgdma_0_dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (msgdma_0_dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (msgdma_0_dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (msgdma_0_dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (msgdma_0_dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (msgdma_0_dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (msgdma_0_dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (msgdma_0_dma_write_master_burstcount),                                         //                          .burstcount
		.av_byteenable         (msgdma_0_dma_write_master_byteenable),                                         //                          .byteenable
		.av_write              (msgdma_0_dma_write_master_write),                                              //                          .write
		.av_writedata          (msgdma_0_dma_write_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (11),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (14),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_if_lpddr2_emif_0_avl_translator (
		.clk                   (mem_if_lpddr2_emif_0_afi_clk_clk),                                                    //                      clk.clk
		.reset                 (rst_controller_006_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount         (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (~mem_if_lpddr2_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) master_0_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_50_clk),                                                                  //       clk.clk
		.reset            (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.av_address       (master_0_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (master_0_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (master_0_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (master_0_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (master_0_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (master_0_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (master_0_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (master_0_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (master_0_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (master_0_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (master_0_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                        //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                        //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_50_clk),                                                                                       //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.av_address       (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (mux_pipeline_007_source0_valid),                                                                   //        rp.valid
		.rp_data          (mux_pipeline_007_source0_data),                                                                    //          .data
		.rp_channel       (mux_pipeline_007_source0_channel),                                                                 //          .channel
		.rp_startofpacket (mux_pipeline_007_source0_startofpacket),                                                           //          .startofpacket
		.rp_endofpacket   (mux_pipeline_007_source0_endofpacket),                                                             //          .endofpacket
		.rp_ready         (mux_pipeline_007_source0_ready)                                                                    //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_source0_ready),                                                                    //              cp.ready
		.cp_valid                (agent_pipeline_source0_valid),                                                                    //                .valid
		.cp_data                 (agent_pipeline_source0_data),                                                                     //                .data
		.cp_startofpacket        (agent_pipeline_source0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (agent_pipeline_source0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (agent_pipeline_source0_channel),                                                                  //                .channel
		.rf_sink_ready           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_002_source0_ready),                                                                   //              cp.ready
		.cp_valid                (agent_pipeline_002_source0_valid),                                                                   //                .valid
		.cp_data                 (agent_pipeline_002_source0_data),                                                                    //                .data
		.cp_startofpacket        (agent_pipeline_002_source0_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (agent_pipeline_002_source0_endofpacket),                                                             //                .endofpacket
		.cp_channel              (agent_pipeline_002_source0_channel),                                                                 //                .channel
		.rf_sink_ready           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_lpddr2_emif_0_afi_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_004_source0_ready),                                                            //              cp.ready
		.cp_valid                (agent_pipeline_004_source0_valid),                                                            //                .valid
		.cp_data                 (agent_pipeline_004_source0_data),                                                             //                .data
		.cp_startofpacket        (agent_pipeline_004_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (agent_pipeline_004_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (agent_pipeline_004_source0_channel),                                                          //                .channel
		.rf_sink_ready           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),                                                      //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (152),
		.PKT_PROTECTION_L          (150),
		.PKT_BEGIN_BURST           (145),
		.PKT_BURSTWRAP_H           (137),
		.PKT_BURSTWRAP_L           (124),
		.PKT_BURST_SIZE_H          (140),
		.PKT_BURST_SIZE_L          (138),
		.PKT_BURST_TYPE_H          (142),
		.PKT_BURST_TYPE_L          (141),
		.PKT_BYTE_CNT_H            (123),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (147),
		.PKT_SRC_ID_L              (147),
		.PKT_DEST_ID_H             (148),
		.PKT_DEST_ID_L             (148),
		.PKT_THREAD_ID_H           (149),
		.PKT_THREAD_ID_L           (149),
		.PKT_CACHE_H               (156),
		.PKT_CACHE_L               (153),
		.PKT_DATA_SIDEBAND_H       (144),
		.PKT_DATA_SIDEBAND_L       (144),
		.PKT_QOS_H                 (146),
		.PKT_QOS_L                 (146),
		.PKT_ADDR_SIDEBAND_H       (143),
		.PKT_ADDR_SIDEBAND_L       (143),
		.ST_DATA_W                 (159),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (9),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (16383),
		.CACHE_VALUE               (4'b0000)
	) msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent (
		.clk              (mem_if_lpddr2_emif_0_afi_clk_clk),                                                     //       clk.clk
		.reset            (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (msgdma_0_dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (msgdma_0_dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (msgdma_0_dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (msgdma_0_dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (msgdma_0_dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (msgdma_0_dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (msgdma_0_dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (msgdma_0_dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (msgdma_0_dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (mux_pipeline_010_source0_valid),                                                       //        rp.valid
		.rp_data          (mux_pipeline_010_source0_data),                                                        //          .data
		.rp_channel       (mux_pipeline_010_source0_channel),                                                     //          .channel
		.rp_startofpacket (mux_pipeline_010_source0_startofpacket),                                               //          .startofpacket
		.rp_endofpacket   (mux_pipeline_010_source0_endofpacket),                                                 //          .endofpacket
		.rp_ready         (mux_pipeline_010_source0_ready)                                                        //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (152),
		.PKT_PROTECTION_L          (150),
		.PKT_BEGIN_BURST           (145),
		.PKT_BURSTWRAP_H           (137),
		.PKT_BURSTWRAP_L           (124),
		.PKT_BURST_SIZE_H          (140),
		.PKT_BURST_SIZE_L          (138),
		.PKT_BURST_TYPE_H          (142),
		.PKT_BURST_TYPE_L          (141),
		.PKT_BYTE_CNT_H            (123),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (147),
		.PKT_SRC_ID_L              (147),
		.PKT_DEST_ID_H             (148),
		.PKT_DEST_ID_L             (148),
		.PKT_THREAD_ID_H           (149),
		.PKT_THREAD_ID_L           (149),
		.PKT_CACHE_H               (156),
		.PKT_CACHE_L               (153),
		.PKT_DATA_SIDEBAND_H       (144),
		.PKT_DATA_SIDEBAND_L       (144),
		.PKT_QOS_H                 (146),
		.PKT_QOS_L                 (146),
		.PKT_ADDR_SIDEBAND_H       (143),
		.PKT_ADDR_SIDEBAND_L       (143),
		.ST_DATA_W                 (159),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (9),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (16383),
		.CACHE_VALUE               (4'b0000)
	) msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent (
		.clk              (mem_if_lpddr2_emif_0_afi_clk_clk),                                                      //       clk.clk
		.reset            (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (msgdma_0_dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (msgdma_0_dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (msgdma_0_dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (msgdma_0_dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (msgdma_0_dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (msgdma_0_dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (msgdma_0_dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (msgdma_0_dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (msgdma_0_dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (mux_pipeline_011_source0_valid),                                                        //        rp.valid
		.rp_data          (mux_pipeline_011_source0_data),                                                         //          .data
		.rp_channel       (mux_pipeline_011_source0_channel),                                                      //          .channel
		.rp_startofpacket (mux_pipeline_011_source0_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (mux_pipeline_011_source0_endofpacket),                                                  //          .endofpacket
		.rp_ready         (mux_pipeline_011_source0_ready)                                                         //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (145),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (147),
		.PKT_SRC_ID_L              (147),
		.PKT_DEST_ID_H             (148),
		.PKT_DEST_ID_L             (148),
		.PKT_BURSTWRAP_H           (137),
		.PKT_BURSTWRAP_L           (124),
		.PKT_BYTE_CNT_H            (123),
		.PKT_BYTE_CNT_L            (110),
		.PKT_PROTECTION_H          (152),
		.PKT_PROTECTION_L          (150),
		.PKT_RESPONSE_STATUS_H     (158),
		.PKT_RESPONSE_STATUS_L     (157),
		.PKT_BURST_SIZE_H          (140),
		.PKT_BURST_SIZE_L          (138),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (159),
		.AVS_BURSTCOUNT_W          (14),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_lpddr2_emif_0_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_006_source0_ready),                                                              //              cp.ready
		.cp_valid                (agent_pipeline_006_source0_valid),                                                              //                .valid
		.cp_data                 (agent_pipeline_006_source0_data),                                                               //                .data
		.cp_startofpacket        (agent_pipeline_006_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_006_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (agent_pipeline_006_source0_channel),                                                            //                .channel
		.rf_sink_ready           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (160),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	q_sys_addr_router addr_router (
		.sink_ready         (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk),                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	q_sys_addr_router_001 addr_router_001 (
		.sink_ready         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (master_driver_msgdma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk),                                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                        //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                        //          .valid
		.src_data           (addr_router_001_src_data),                                                                         //          .data
		.src_channel        (addr_router_001_src_channel),                                                                      //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                                   //          .endofpacket
	);

	q_sys_id_router id_router (
		.sink_ready         (agent_pipeline_001_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_001_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_001_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_001_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_001_source0_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_src_ready),                      //       src.ready
		.src_valid          (id_router_src_valid),                      //          .valid
		.src_data           (id_router_src_data),                       //          .data
		.src_channel        (id_router_src_channel),                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                 //          .endofpacket
	);

	q_sys_id_router id_router_001 (
		.sink_ready         (agent_pipeline_003_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_003_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_003_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_003_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_003_source0_endofpacket),   //          .endofpacket
		.clk                (clk_50_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                  //       src.ready
		.src_valid          (id_router_001_src_valid),                  //          .valid
		.src_data           (id_router_001_src_data),                   //          .data
		.src_channel        (id_router_001_src_channel),                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)             //          .endofpacket
	);

	q_sys_id_router_002 id_router_002 (
		.sink_ready         (agent_pipeline_005_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_005_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_005_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_005_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_005_source0_endofpacket),   //          .endofpacket
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),         //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                  //       src.ready
		.src_valid          (id_router_002_src_valid),                  //          .valid
		.src_data           (id_router_002_src_data),                   //          .data
		.src_channel        (id_router_002_src_channel),                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)             //          .endofpacket
	);

	q_sys_addr_router_002 addr_router_002 (
		.sink_ready         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (msgdma_0_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	q_sys_addr_router_002 addr_router_003 (
		.sink_ready         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (msgdma_0_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	q_sys_id_router_003 id_router_003 (
		.sink_ready         (agent_pipeline_007_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_007_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_007_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_007_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_007_source0_endofpacket),   //          .endofpacket
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),         //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                  //       src.ready
		.src_valid          (id_router_003_src_valid),                  //          .valid
		.src_data           (id_router_003_src_data),                   //          .data
		.src_channel        (id_router_003_src_channel),                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)             //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (20),
		.PIPELINED                 (0),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (3),
		.VALID_WIDTH               (1),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_50_clk),                                 //       clk.clk
		.reset                  (rst_controller_002_reset_out_reset),         // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),                      //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),                      //          .valid
		.cmd_sink_data          (addr_router_src_data),                       //          .data
		.cmd_sink_channel       (addr_router_src_channel),                    //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),              //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),                //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),                      //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),                       //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),                    //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),              //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),                //          .endofpacket
		.cmd_src_valid          (limiter_cmd_src_valid),                      //          .valid
		.rsp_sink_ready         (limiter_pipeline_001_source0_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.rsp_sink_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.rsp_sink_data          (limiter_pipeline_001_source0_data),          //          .data
		.rsp_sink_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),                      //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),                      //          .valid
		.rsp_src_data           (limiter_rsp_src_data),                       //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),                    //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),              //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket)                 //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (master_driver_msgdma_0_reset_source_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                            // reset_in1.reset
		.reset_in2  (~mem_if_lpddr2_emif_0_afi_reset_reset),     // reset_in2.reset
		.clk        (),                                          //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),            // reset_out.reset
		.reset_in3  (1'b0),                                      // (terminated)
		.reset_in4  (1'b0),                                      // (terminated)
		.reset_in5  (1'b0),                                      // (terminated)
		.reset_in6  (1'b0),                                      // (terminated)
		.reset_in7  (1'b0),                                      // (terminated)
		.reset_in8  (1'b0),                                      // (terminated)
		.reset_in9  (1'b0),                                      // (terminated)
		.reset_in10 (1'b0),                                      // (terminated)
		.reset_in11 (1'b0),                                      // (terminated)
		.reset_in12 (1'b0),                                      // (terminated)
		.reset_in13 (1'b0),                                      // (terminated)
		.reset_in14 (1'b0),                                      // (terminated)
		.reset_in15 (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_50_reset_n),                     // reset_in0.reset
		.reset_in1  (~mem_if_lpddr2_emif_0_afi_reset_reset), // reset_in1.reset
		.clk        (),                                      //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_50_reset_n),                  // reset_in0.reset
		.clk        (clk_50_clk),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_50_reset_n),                     // reset_in0.reset
		.reset_in1  (~mem_if_lpddr2_emif_0_afi_reset_reset), // reset_in1.reset
		.clk        (clk_50_clk),                            //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (master_driver_msgdma_0_reset_source_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                            // reset_in1.reset
		.reset_in2  (~mem_if_lpddr2_emif_0_afi_reset_reset),     // reset_in2.reset
		.clk        (mem_if_lpddr2_emif_0_afi_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),        // reset_out.reset
		.reset_in3  (1'b0),                                      // (terminated)
		.reset_in4  (1'b0),                                      // (terminated)
		.reset_in5  (1'b0),                                      // (terminated)
		.reset_in6  (1'b0),                                      // (terminated)
		.reset_in7  (1'b0),                                      // (terminated)
		.reset_in8  (1'b0),                                      // (terminated)
		.reset_in9  (1'b0),                                      // (terminated)
		.reset_in10 (1'b0),                                      // (terminated)
		.reset_in11 (1'b0),                                      // (terminated)
		.reset_in12 (1'b0),                                      // (terminated)
		.reset_in13 (1'b0),                                      // (terminated)
		.reset_in14 (1'b0),                                      // (terminated)
		.reset_in15 (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_006 (
		.reset_in0  (~mem_if_lpddr2_emif_0_afi_reset_reset), // reset_in0.reset
		.clk        (mem_if_lpddr2_emif_0_afi_clk_clk),      //       clk.clk
		.reset_out  (rst_controller_006_reset_out_reset),    // reset_out.reset
		.reset_in1  (1'b0),                                  // (terminated)
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	q_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_50_clk),                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.sink_ready         (limiter_pipeline_source0_ready),         //      sink.ready
		.sink_channel       (limiter_pipeline_source0_channel),       //          .channel
		.sink_data          (limiter_pipeline_source0_data),          //          .data
		.sink_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.sink_valid         (limiter_pipeline_source0_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),              //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),               //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),        //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),              //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),              //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),               //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),            //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),        //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),              //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),              //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),               //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),            //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),      //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)         //          .endofpacket
	);

	q_sys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_50_clk),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	q_sys_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (mem_if_lpddr2_emif_0_afi_clk_clk),       //       clk.clk
		.reset               (rst_controller_005_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),       //          .endofpacket
		.sink0_ready         (mux_pipeline_002_source0_ready),         //     sink0.ready
		.sink0_valid         (mux_pipeline_002_source0_valid),         //          .valid
		.sink0_channel       (mux_pipeline_002_source0_channel),       //          .channel
		.sink0_data          (mux_pipeline_002_source0_data),          //          .data
		.sink0_startofpacket (mux_pipeline_002_source0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_002_source0_endofpacket),   //          .endofpacket
		.sink1_ready         (mux_pipeline_003_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_003_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_003_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_003_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_003_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_003_source0_endofpacket)    //          .endofpacket
	);

	q_sys_cmd_xbar_demux_001 rsp_xbar_demux (
		.clk                (clk_50_clk),                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	q_sys_cmd_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_50_clk),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	q_sys_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	q_sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_50_clk),                             //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                 //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                 //          .valid
		.src_data            (rsp_xbar_mux_src_data),                  //          .data
		.src_channel         (rsp_xbar_mux_src_channel),               //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),         //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),           //          .endofpacket
		.sink0_ready         (mux_pipeline_004_source0_ready),         //     sink0.ready
		.sink0_valid         (mux_pipeline_004_source0_valid),         //          .valid
		.sink0_channel       (mux_pipeline_004_source0_channel),       //          .channel
		.sink0_data          (mux_pipeline_004_source0_data),          //          .data
		.sink0_startofpacket (mux_pipeline_004_source0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_004_source0_endofpacket),   //          .endofpacket
		.sink1_ready         (mux_pipeline_005_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_005_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_005_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_005_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_005_source0_endofpacket),   //          .endofpacket
		.sink2_ready         (mux_pipeline_006_source0_ready),         //     sink2.ready
		.sink2_valid         (mux_pipeline_006_source0_valid),         //          .valid
		.sink2_channel       (mux_pipeline_006_source0_channel),       //          .channel
		.sink2_data          (mux_pipeline_006_source0_data),          //          .data
		.sink2_startofpacket (mux_pipeline_006_source0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (mux_pipeline_006_source0_endofpacket)    //          .endofpacket
	);

	q_sys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	q_sys_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	q_sys_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (mem_if_lpddr2_emif_0_afi_clk_clk),       //       clk.clk
		.reset               (rst_controller_006_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),       //          .endofpacket
		.sink0_ready         (mux_pipeline_008_source0_ready),         //     sink0.ready
		.sink0_valid         (mux_pipeline_008_source0_valid),         //          .valid
		.sink0_channel       (mux_pipeline_008_source0_channel),       //          .channel
		.sink0_data          (mux_pipeline_008_source0_data),          //          .data
		.sink0_startofpacket (mux_pipeline_008_source0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_008_source0_endofpacket),   //          .endofpacket
		.sink1_ready         (mux_pipeline_009_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_009_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_009_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_009_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_009_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_009_source0_endofpacket)    //          .endofpacket
	);

	q_sys_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (mem_if_lpddr2_emif_0_afi_clk_clk),      //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (3),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_50_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (mem_if_lpddr2_emif_0_afi_clk_clk),   //       out_clk.clk
		.out_reset         (rst_controller_005_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src2_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src2_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src2_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src2_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (3),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_50_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_lpddr2_emif_0_afi_clk_clk),      //       out_clk.clk
		.out_reset         (rst_controller_005_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (3),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (mem_if_lpddr2_emif_0_afi_clk_clk),      //        in_clk.clk
		.in_reset          (rst_controller_005_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_50_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_002_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_002_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_002_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_002_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (3),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (mem_if_lpddr2_emif_0_afi_clk_clk),      //        in_clk.clk
		.in_reset          (rst_controller_005_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_50_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_002_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_002_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_002_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_002_src1_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),     // cr0_reset.reset
		.in_ready          (limiter_cmd_src_ready),                  //     sink0.ready
		.in_valid          (limiter_cmd_src_valid),                  //          .valid
		.in_startofpacket  (limiter_cmd_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (limiter_cmd_src_endofpacket),            //          .endofpacket
		.in_data           (limiter_cmd_src_data),                   //          .data
		.in_channel        (limiter_cmd_src_channel),                //          .channel
		.out_ready         (limiter_pipeline_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_source0_data),          //          .data
		.out_channel       (limiter_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_001 (
		.clk               (clk_50_clk),                                 //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_mux_src_ready),                     //     sink0.ready
		.in_valid          (rsp_xbar_mux_src_valid),                     //          .valid
		.in_startofpacket  (rsp_xbar_mux_src_startofpacket),             //          .startofpacket
		.in_endofpacket    (rsp_xbar_mux_src_endofpacket),               //          .endofpacket
		.in_data           (rsp_xbar_mux_src_data),                      //          .data
		.in_channel        (rsp_xbar_mux_src_channel),                   //          .channel
		.out_ready         (limiter_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_001_source0_data),          //          .data
		.out_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline (
		.clk               (clk_50_clk),                           //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),   // cr0_reset.reset
		.in_ready          (mux_pipeline_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_source0_data),            //          .data
		.in_channel        (mux_pipeline_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_source0_data),          //          .data
		.out_channel       (agent_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.out_error         (),                                     // (terminated)
		.in_error          (1'b0)                                  // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_001 (
		.clk               (clk_50_clk),                                                                            //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),                                                    // cr0_reset.reset
		.in_ready          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (master_driver_msgdma_0_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_001_source0_ready),                                                      //   source0.ready
		.out_valid         (agent_pipeline_001_source0_valid),                                                      //          .valid
		.out_startofpacket (agent_pipeline_001_source0_startofpacket),                                              //          .startofpacket
		.out_endofpacket   (agent_pipeline_001_source0_endofpacket),                                                //          .endofpacket
		.out_data          (agent_pipeline_001_source0_data),                                                       //          .data
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_channel       (),                                                                                      // (terminated)
		.in_channel        (1'b0)                                                                                   // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_002 (
		.clk               (clk_50_clk),                               //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),       // cr0_reset.reset
		.in_ready          (mux_pipeline_001_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_001_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_001_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_001_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_001_source0_data),            //          .data
		.in_channel        (mux_pipeline_001_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_002_source0_data),          //          .data
		.out_channel       (agent_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_003 (
		.clk               (clk_50_clk),                                                                               //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),                                                       // cr0_reset.reset
		.in_ready          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (product_info_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_003_source0_ready),                                                         //   source0.ready
		.out_valid         (agent_pipeline_003_source0_valid),                                                         //          .valid
		.out_startofpacket (agent_pipeline_003_source0_startofpacket),                                                 //          .startofpacket
		.out_endofpacket   (agent_pipeline_003_source0_endofpacket),                                                   //          .endofpacket
		.out_data          (agent_pipeline_003_source0_data),                                                          //          .data
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_channel       (),                                                                                         // (terminated)
		.in_channel        (1'b0)                                                                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_004 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),         //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),       // cr0_reset.reset
		.in_ready          (cmd_xbar_mux_002_src_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_mux_002_src_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_mux_002_src_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_002_src_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_mux_002_src_data),                //          .data
		.in_channel        (cmd_xbar_mux_002_src_channel),             //          .channel
		.out_ready         (agent_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_004_source0_data),          //          .data
		.out_channel       (agent_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_005 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),                                                  //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),                                                // cr0_reset.reset
		.in_ready          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (msgdma_0_mm_bridge_slv_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_005_source0_ready),                                                  //   source0.ready
		.out_valid         (agent_pipeline_005_source0_valid),                                                  //          .valid
		.out_startofpacket (agent_pipeline_005_source0_startofpacket),                                          //          .startofpacket
		.out_endofpacket   (agent_pipeline_005_source0_endofpacket),                                            //          .endofpacket
		.out_data          (agent_pipeline_005_source0_data),                                                   //          .data
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_channel       (),                                                                                  // (terminated)
		.in_channel        (1'b0)                                                                               // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_006 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),         //       cr0.clk
		.reset             (rst_controller_006_reset_out_reset),       // cr0_reset.reset
		.in_ready          (cmd_xbar_mux_003_src_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_mux_003_src_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_mux_003_src_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_003_src_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_mux_003_src_data),                //          .data
		.in_channel        (cmd_xbar_mux_003_src_channel),             //          .channel
		.out_ready         (agent_pipeline_006_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_006_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_006_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_006_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_006_source0_data),          //          .data
		.out_channel       (agent_pipeline_006_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_007 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),                                                    //       cr0.clk
		.reset             (rst_controller_006_reset_out_reset),                                                  // cr0_reset.reset
		.in_ready          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (mem_if_lpddr2_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_007_source0_ready),                                                    //   source0.ready
		.out_valid         (agent_pipeline_007_source0_valid),                                                    //          .valid
		.out_startofpacket (agent_pipeline_007_source0_startofpacket),                                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_007_source0_endofpacket),                                              //          .endofpacket
		.out_data          (agent_pipeline_007_source0_data),                                                     //          .data
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_channel       (),                                                                                    // (terminated)
		.in_channel        (1'b0)                                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline (
		.clk               (clk_50_clk),                         //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset), // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_src0_data),           //          .data
		.in_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_source0_data),          //          .data
		.out_channel       (mux_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                               // (terminated)
		.out_empty         (),                                   // (terminated)
		.out_error         (),                                   // (terminated)
		.in_error          (1'b0)                                // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_001 (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),     // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src1_ready),              //     sink0.ready
		.in_valid          (cmd_xbar_demux_src1_valid),              //          .valid
		.in_startofpacket  (cmd_xbar_demux_src1_startofpacket),      //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src1_endofpacket),        //          .endofpacket
		.in_data           (cmd_xbar_demux_src1_data),               //          .data
		.in_channel        (cmd_xbar_demux_src1_channel),            //          .channel
		.out_ready         (mux_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_001_source0_data),          //          .data
		.out_channel       (mux_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_002 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_out_ready),                      //     sink0.ready
		.in_valid          (crosser_out_valid),                      //          .valid
		.in_startofpacket  (crosser_out_startofpacket),              //          .startofpacket
		.in_endofpacket    (crosser_out_endofpacket),                //          .endofpacket
		.in_data           (crosser_out_data),                       //          .data
		.in_channel        (crosser_out_channel),                    //          .channel
		.out_ready         (mux_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_002_source0_data),          //          .data
		.out_channel       (mux_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_003 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_001_out_ready),                  //     sink0.ready
		.in_valid          (crosser_001_out_valid),                  //          .valid
		.in_startofpacket  (crosser_001_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_001_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_001_out_data),                   //          .data
		.in_channel        (crosser_001_out_channel),                //          .channel
		.out_ready         (mux_pipeline_003_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_003_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_003_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_003_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_003_source0_data),          //          .data
		.out_channel       (mux_pipeline_003_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_004 (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),     // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),              //     sink0.ready
		.in_valid          (rsp_xbar_demux_src0_valid),              //          .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),        //          .endofpacket
		.in_data           (rsp_xbar_demux_src0_data),               //          .data
		.in_channel        (rsp_xbar_demux_src0_channel),            //          .channel
		.out_ready         (mux_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_004_source0_data),          //          .data
		.out_channel       (mux_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_005 (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),     // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_001_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_001_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_001_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_001_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_005_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_005_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_005_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_005_source0_data),          //          .data
		.out_channel       (mux_pipeline_005_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_006 (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_002_out_ready),                  //     sink0.ready
		.in_valid          (crosser_002_out_valid),                  //          .valid
		.in_startofpacket  (crosser_002_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_002_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_002_out_data),                   //          .data
		.in_channel        (crosser_002_out_channel),                //          .channel
		.out_ready         (mux_pipeline_006_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_006_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_006_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_006_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_006_source0_data),          //          .data
		.out_channel       (mux_pipeline_006_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (103),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (3),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_007 (
		.clk               (clk_50_clk),                             //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),     // cr0_reset.reset
		.in_ready          (crosser_003_out_ready),                  //     sink0.ready
		.in_valid          (crosser_003_out_valid),                  //          .valid
		.in_startofpacket  (crosser_003_out_startofpacket),          //          .startofpacket
		.in_endofpacket    (crosser_003_out_endofpacket),            //          .endofpacket
		.in_data           (crosser_003_out_data),                   //          .data
		.in_channel        (crosser_003_out_channel),                //          .channel
		.out_ready         (mux_pipeline_007_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_007_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_007_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_007_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_007_source0_data),          //          .data
		.out_channel       (mux_pipeline_007_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_008 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_006_reset_out_reset),     // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_002_src0_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_002_src0_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_002_src0_data),           //          .data
		.in_channel        (cmd_xbar_demux_002_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_008_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_008_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_008_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_008_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_008_source0_data),          //          .data
		.out_channel       (mux_pipeline_008_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_009 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_006_reset_out_reset),     // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_003_src0_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_003_src0_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_003_src0_data),           //          .data
		.in_channel        (cmd_xbar_demux_003_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_009_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_009_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_009_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_009_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_009_source0_data),          //          .data
		.out_channel       (mux_pipeline_009_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_010 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),     // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_003_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_003_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_003_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_003_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_010_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_010_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_010_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_010_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_010_source0_data),          //          .data
		.out_channel       (mux_pipeline_010_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (159),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_011 (
		.clk               (mem_if_lpddr2_emif_0_afi_clk_clk),       //       cr0.clk
		.reset             (rst_controller_005_reset_out_reset),     // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_003_src1_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_003_src1_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_003_src1_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_003_src1_data),           //          .data
		.in_channel        (rsp_xbar_demux_003_src1_channel),        //          .channel
		.out_ready         (mux_pipeline_011_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_011_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_011_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_011_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_011_source0_data),          //          .data
		.out_channel       (mux_pipeline_011_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	q_sys_irq_mapper irq_mapper (
		.clk           (clk_50_clk),                                    //       clk.clk
		.reset         (rst_controller_003_reset_out_reset),            // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),                      // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),                      // receiver1.irq
		.sender_irq    (master_driver_msgdma_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (mem_if_lpddr2_emif_0_afi_clk_clk),   //       receiver_clk.clk
		.sender_clk     (clk_50_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (mem_if_lpddr2_emif_0_afi_clk_clk),   //       receiver_clk.clk
		.sender_clk     (clk_50_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

endmodule
